--------------------------------------------------------------------------------
--                         ModuloCounter_16_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_16_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of ModuloCounter_16_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(3 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 15 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1589838
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1589838 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1589838 is
signal XX_m1589839 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m1589839 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m1589839 <= X ;
   YY_m1589839 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid1589842
--                   (IntAdderClassical_33_f500_uid1589844)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid1589842 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid1589842 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1589838 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid1589842 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1589838  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
   RoundingAdder: IntAdder_33_f500_uid1589842  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound   ,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_16_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_16_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_16_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
         iS_11 when "1011",
         iS_12 when "1100",
         iS_13 when "1101",
         iS_14 when "1110",
         iS_15 when "1111",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_5_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_5_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_5_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid1590613_RightShifter
--                (RightShifter_24_by_max_26_F250_uid1590615)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1590613_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1590613_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid1590618
--                  (IntAdderAlternative_27_f250_uid1590622)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid1590618 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid1590618 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid1590625
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid1590625 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid1590625 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid1590628
--                   (IntAdderClassical_34_f250_uid1590630)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid1590628 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid1590628 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid1590613
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1590613 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1590613 is
   component FPAdd_8_23_uid1590613_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid1590618 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid1590625 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid1590628 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid1590613_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid1590618  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid1590625  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid1590628  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid1590613 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid1590613  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_11_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_11_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_11_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_10_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_10_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_10_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_9_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_9_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_9_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid1591691_RightShifter
--                (RightShifter_24_by_max_26_F250_uid1591693)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1591691_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1591691_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid1591696
--                  (IntAdderAlternative_27_f250_uid1591700)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid1591696 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid1591696 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid1591703
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid1591703 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid1591703 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid1591706
--                   (IntAdderClassical_34_f250_uid1591708)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid1591706 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid1591706 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid1591691
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1591691 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1591691 is
   component FPAdd_8_23_uid1591691_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid1591696 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid1591703 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid1591706 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid1591691_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid1591696  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid1591703  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid1591706  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid1591691 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid1591691  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_12_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_12_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_12_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
         iS_11 when "1011",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                            SelFunctionTable_r8
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity SelFunctionTable_r8 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(6 downto 0);
          Y : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of SelFunctionTable_r8 is
begin
  with X select  Y <= 
   "0000" when "0000000",
   "0000" when "0000001",
   "0000" when "0000010",
   "0000" when "0000011",
   "0001" when "0000100",
   "0001" when "0000101",
   "0001" when "0000110",
   "0001" when "0000111",
   "0001" when "0001000",
   "0001" when "0001001",
   "0001" when "0001010",
   "0001" when "0001011",
   "0010" when "0001100",
   "0010" when "0001101",
   "0010" when "0001110",
   "0010" when "0001111",
   "0011" when "0010000",
   "0011" when "0010001",
   "0010" when "0010010",
   "0010" when "0010011",
   "0011" when "0010100",
   "0011" when "0010101",
   "0011" when "0010110",
   "0011" when "0010111",
   "0100" when "0011000",
   "0100" when "0011001",
   "0011" when "0011010",
   "0011" when "0011011",
   "0101" when "0011100",
   "0100" when "0011101",
   "0100" when "0011110",
   "0100" when "0011111",
   "0101" when "0100000",
   "0101" when "0100001",
   "0101" when "0100010",
   "0100" when "0100011",
   "0110" when "0100100",
   "0110" when "0100101",
   "0101" when "0100110",
   "0101" when "0100111",
   "0111" when "0101000",
   "0110" when "0101001",
   "0110" when "0101010",
   "0101" when "0101011",
   "0111" when "0101100",
   "0111" when "0101101",
   "0110" when "0101110",
   "0110" when "0101111",
   "0111" when "0110000",
   "0111" when "0110001",
   "0111" when "0110010",
   "0110" when "0110011",
   "0111" when "0110100",
   "0111" when "0110101",
   "0111" when "0110110",
   "0111" when "0110111",
   "0111" when "0111000",
   "0111" when "0111001",
   "0111" when "0111010",
   "0111" when "0111011",
   "0111" when "0111100",
   "0111" when "0111101",
   "0111" when "0111110",
   "0111" when "0111111",
   "1001" when "1000000",
   "1001" when "1000001",
   "1001" when "1000010",
   "1001" when "1000011",
   "1001" when "1000100",
   "1001" when "1000101",
   "1001" when "1000110",
   "1001" when "1000111",
   "1001" when "1001000",
   "1001" when "1001001",
   "1001" when "1001010",
   "1001" when "1001011",
   "1001" when "1001100",
   "1001" when "1001101",
   "1001" when "1001110",
   "1001" when "1001111",
   "1001" when "1010000",
   "1001" when "1010001",
   "1010" when "1010010",
   "1010" when "1010011",
   "1001" when "1010100",
   "1010" when "1010101",
   "1010" when "1010110",
   "1010" when "1010111",
   "1010" when "1011000",
   "1010" when "1011001",
   "1011" when "1011010",
   "1011" when "1011011",
   "1011" when "1011100",
   "1011" when "1011101",
   "1011" when "1011110",
   "1011" when "1011111",
   "1011" when "1100000",
   "1011" when "1100001",
   "1100" when "1100010",
   "1100" when "1100011",
   "1100" when "1100100",
   "1100" when "1100101",
   "1100" when "1100110",
   "1100" when "1100111",
   "1100" when "1101000",
   "1101" when "1101001",
   "1101" when "1101010",
   "1101" when "1101011",
   "1101" when "1101100",
   "1101" when "1101101",
   "1101" when "1101110",
   "1101" when "1101111",
   "1110" when "1110000",
   "1110" when "1110001",
   "1110" when "1110010",
   "1110" when "1110011",
   "1110" when "1110100",
   "1110" when "1110101",
   "1110" when "1110110",
   "1110" when "1110111",
   "1111" when "1111000",
   "1111" when "1111001",
   "1111" when "1111010",
   "1111" when "1111011",
   "1111" when "1111100",
   "1111" when "1111101",
   "1111" when "1111110",
   "1111" when "1111111",
   "----" when others;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
   component SelFunctionTable_r8 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(6 downto 0);
             Y : out std_logic_vector(3 downto 0)   );
   end component;

signal partialFX : std_logic_vector(23 downto 0) := (others => '0');
signal partialFY : std_logic_vector(23 downto 0) := (others => '0');
signal expR0, expR0_d1, expR0_d2, expR0_d3, expR0_d4, expR0_d5, expR0_d6, expR0_d7, expR0_d8, expR0_d9, expR0_d10, expR0_d11 : std_logic_vector(9 downto 0) := (others => '0');
signal sR, sR_d1, sR_d2, sR_d3, sR_d4, sR_d5, sR_d6, sR_d7, sR_d8, sR_d9, sR_d10, sR_d11, sR_d12 : std_logic := '0';
signal exnXY : std_logic_vector(3 downto 0) := (others => '0');
signal exnR0, exnR0_d1, exnR0_d2, exnR0_d3, exnR0_d4, exnR0_d5, exnR0_d6, exnR0_d7, exnR0_d8, exnR0_d9, exnR0_d10, exnR0_d11, exnR0_d12 : std_logic_vector(1 downto 0) := (others => '0');
signal fY, fY_d1, fY_d2, fY_d3, fY_d4, fY_d5, fY_d6, fY_d7, fY_d8, fY_d9 : std_logic_vector(25 downto 0) := (others => '0');
signal fX : std_logic_vector(26 downto 0) := (others => '0');
signal w9, w9_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel9 : std_logic_vector(6 downto 0) := (others => '0');
signal q9, q9_d1, q9_d2, q9_d3, q9_d4, q9_d5, q9_d6, q9_d7, q9_d8, q9_d9 : std_logic_vector(3 downto 0) := (others => '0');
signal w9pad : std_logic_vector(29 downto 0) := (others => '0');
signal w8fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec8 : std_logic_vector(29 downto 0) := (others => '0');
signal w8full : std_logic_vector(29 downto 0) := (others => '0');
signal w8, w8_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel8 : std_logic_vector(6 downto 0) := (others => '0');
signal q8, q8_d1, q8_d2, q8_d3, q8_d4, q8_d5, q8_d6, q8_d7, q8_d8 : std_logic_vector(3 downto 0) := (others => '0');
signal w8pad : std_logic_vector(29 downto 0) := (others => '0');
signal w7fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec7 : std_logic_vector(29 downto 0) := (others => '0');
signal w7full : std_logic_vector(29 downto 0) := (others => '0');
signal w7, w7_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel7 : std_logic_vector(6 downto 0) := (others => '0');
signal q7, q7_d1, q7_d2, q7_d3, q7_d4, q7_d5, q7_d6, q7_d7 : std_logic_vector(3 downto 0) := (others => '0');
signal w7pad : std_logic_vector(29 downto 0) := (others => '0');
signal w6fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec6 : std_logic_vector(29 downto 0) := (others => '0');
signal w6full : std_logic_vector(29 downto 0) := (others => '0');
signal w6, w6_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel6 : std_logic_vector(6 downto 0) := (others => '0');
signal q6, q6_d1, q6_d2, q6_d3, q6_d4, q6_d5, q6_d6 : std_logic_vector(3 downto 0) := (others => '0');
signal w6pad : std_logic_vector(29 downto 0) := (others => '0');
signal w5fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec5 : std_logic_vector(29 downto 0) := (others => '0');
signal w5full : std_logic_vector(29 downto 0) := (others => '0');
signal w5, w5_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel5 : std_logic_vector(6 downto 0) := (others => '0');
signal q5, q5_d1, q5_d2, q5_d3, q5_d4, q5_d5 : std_logic_vector(3 downto 0) := (others => '0');
signal w5pad : std_logic_vector(29 downto 0) := (others => '0');
signal w4fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec4 : std_logic_vector(29 downto 0) := (others => '0');
signal w4full : std_logic_vector(29 downto 0) := (others => '0');
signal w4, w4_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel4 : std_logic_vector(6 downto 0) := (others => '0');
signal q4, q4_d1, q4_d2, q4_d3, q4_d4 : std_logic_vector(3 downto 0) := (others => '0');
signal w4pad : std_logic_vector(29 downto 0) := (others => '0');
signal w3fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec3 : std_logic_vector(29 downto 0) := (others => '0');
signal w3full : std_logic_vector(29 downto 0) := (others => '0');
signal w3, w3_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel3 : std_logic_vector(6 downto 0) := (others => '0');
signal q3, q3_d1, q3_d2, q3_d3 : std_logic_vector(3 downto 0) := (others => '0');
signal w3pad : std_logic_vector(29 downto 0) := (others => '0');
signal w2fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec2 : std_logic_vector(29 downto 0) := (others => '0');
signal w2full : std_logic_vector(29 downto 0) := (others => '0');
signal w2, w2_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel2 : std_logic_vector(6 downto 0) := (others => '0');
signal q2, q2_d1, q2_d2 : std_logic_vector(3 downto 0) := (others => '0');
signal w2pad : std_logic_vector(29 downto 0) := (others => '0');
signal w1fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec1 : std_logic_vector(29 downto 0) := (others => '0');
signal w1full : std_logic_vector(29 downto 0) := (others => '0');
signal w1, w1_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel1 : std_logic_vector(6 downto 0) := (others => '0');
signal q1, q1_d1 : std_logic_vector(3 downto 0) := (others => '0');
signal w1pad : std_logic_vector(29 downto 0) := (others => '0');
signal w0fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec0 : std_logic_vector(29 downto 0) := (others => '0');
signal w0full : std_logic_vector(29 downto 0) := (others => '0');
signal w0, w0_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal q0 : std_logic_vector(3 downto 0) := (others => '0');
signal qP9 : std_logic_vector(2 downto 0) := (others => '0');
signal qM9 : std_logic_vector(2 downto 0) := (others => '0');
signal qP8 : std_logic_vector(2 downto 0) := (others => '0');
signal qM8 : std_logic_vector(2 downto 0) := (others => '0');
signal qP7 : std_logic_vector(2 downto 0) := (others => '0');
signal qM7 : std_logic_vector(2 downto 0) := (others => '0');
signal qP6 : std_logic_vector(2 downto 0) := (others => '0');
signal qM6 : std_logic_vector(2 downto 0) := (others => '0');
signal qP5 : std_logic_vector(2 downto 0) := (others => '0');
signal qM5 : std_logic_vector(2 downto 0) := (others => '0');
signal qP4 : std_logic_vector(2 downto 0) := (others => '0');
signal qM4 : std_logic_vector(2 downto 0) := (others => '0');
signal qP3 : std_logic_vector(2 downto 0) := (others => '0');
signal qM3 : std_logic_vector(2 downto 0) := (others => '0');
signal qP2 : std_logic_vector(2 downto 0) := (others => '0');
signal qM2 : std_logic_vector(2 downto 0) := (others => '0');
signal qP1 : std_logic_vector(2 downto 0) := (others => '0');
signal qM1 : std_logic_vector(2 downto 0) := (others => '0');
signal qP0 : std_logic_vector(2 downto 0) := (others => '0');
signal qM0 : std_logic_vector(2 downto 0) := (others => '0');
signal qP : std_logic_vector(29 downto 0) := (others => '0');
signal qM : std_logic_vector(29 downto 0) := (others => '0');
signal fR0, fR0_d1 : std_logic_vector(29 downto 0) := (others => '0');
signal fR : std_logic_vector(28 downto 0) := (others => '0');
signal fRn1, fRn1_d1 : std_logic_vector(26 downto 0) := (others => '0');
signal expR1, expR1_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal round, round_d1 : std_logic := '0';
signal expfrac : std_logic_vector(32 downto 0) := (others => '0');
signal expfracR : std_logic_vector(32 downto 0) := (others => '0');
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
signal exnRfinal : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            expR0_d1 <=  expR0;
            expR0_d2 <=  expR0_d1;
            expR0_d3 <=  expR0_d2;
            expR0_d4 <=  expR0_d3;
            expR0_d5 <=  expR0_d4;
            expR0_d6 <=  expR0_d5;
            expR0_d7 <=  expR0_d6;
            expR0_d8 <=  expR0_d7;
            expR0_d9 <=  expR0_d8;
            expR0_d10 <=  expR0_d9;
            expR0_d11 <=  expR0_d10;
            sR_d1 <=  sR;
            sR_d2 <=  sR_d1;
            sR_d3 <=  sR_d2;
            sR_d4 <=  sR_d3;
            sR_d5 <=  sR_d4;
            sR_d6 <=  sR_d5;
            sR_d7 <=  sR_d6;
            sR_d8 <=  sR_d7;
            sR_d9 <=  sR_d8;
            sR_d10 <=  sR_d9;
            sR_d11 <=  sR_d10;
            sR_d12 <=  sR_d11;
            exnR0_d1 <=  exnR0;
            exnR0_d2 <=  exnR0_d1;
            exnR0_d3 <=  exnR0_d2;
            exnR0_d4 <=  exnR0_d3;
            exnR0_d5 <=  exnR0_d4;
            exnR0_d6 <=  exnR0_d5;
            exnR0_d7 <=  exnR0_d6;
            exnR0_d8 <=  exnR0_d7;
            exnR0_d9 <=  exnR0_d8;
            exnR0_d10 <=  exnR0_d9;
            exnR0_d11 <=  exnR0_d10;
            exnR0_d12 <=  exnR0_d11;
            fY_d1 <=  fY;
            fY_d2 <=  fY_d1;
            fY_d3 <=  fY_d2;
            fY_d4 <=  fY_d3;
            fY_d5 <=  fY_d4;
            fY_d6 <=  fY_d5;
            fY_d7 <=  fY_d6;
            fY_d8 <=  fY_d7;
            fY_d9 <=  fY_d8;
            w9_d1 <=  w9;
            q9_d1 <=  q9;
            q9_d2 <=  q9_d1;
            q9_d3 <=  q9_d2;
            q9_d4 <=  q9_d3;
            q9_d5 <=  q9_d4;
            q9_d6 <=  q9_d5;
            q9_d7 <=  q9_d6;
            q9_d8 <=  q9_d7;
            q9_d9 <=  q9_d8;
            w8_d1 <=  w8;
            q8_d1 <=  q8;
            q8_d2 <=  q8_d1;
            q8_d3 <=  q8_d2;
            q8_d4 <=  q8_d3;
            q8_d5 <=  q8_d4;
            q8_d6 <=  q8_d5;
            q8_d7 <=  q8_d6;
            q8_d8 <=  q8_d7;
            w7_d1 <=  w7;
            q7_d1 <=  q7;
            q7_d2 <=  q7_d1;
            q7_d3 <=  q7_d2;
            q7_d4 <=  q7_d3;
            q7_d5 <=  q7_d4;
            q7_d6 <=  q7_d5;
            q7_d7 <=  q7_d6;
            w6_d1 <=  w6;
            q6_d1 <=  q6;
            q6_d2 <=  q6_d1;
            q6_d3 <=  q6_d2;
            q6_d4 <=  q6_d3;
            q6_d5 <=  q6_d4;
            q6_d6 <=  q6_d5;
            w5_d1 <=  w5;
            q5_d1 <=  q5;
            q5_d2 <=  q5_d1;
            q5_d3 <=  q5_d2;
            q5_d4 <=  q5_d3;
            q5_d5 <=  q5_d4;
            w4_d1 <=  w4;
            q4_d1 <=  q4;
            q4_d2 <=  q4_d1;
            q4_d3 <=  q4_d2;
            q4_d4 <=  q4_d3;
            w3_d1 <=  w3;
            q3_d1 <=  q3;
            q3_d2 <=  q3_d1;
            q3_d3 <=  q3_d2;
            w2_d1 <=  w2;
            q2_d1 <=  q2;
            q2_d2 <=  q2_d1;
            w1_d1 <=  w1;
            q1_d1 <=  q1;
            w0_d1 <=  w0;
            fR0_d1 <=  fR0;
            fRn1_d1 <=  fRn1;
            expR1_d1 <=  expR1;
            round_d1 <=  round;
         end if;
      end process;
   partialFX <= "1" & X(22 downto 0);
   partialFY <= "1" & Y(22 downto 0);
   -- exponent difference, sign and exception combination computed early, to have less bits to pipeline
   expR0 <= ("00" & X(30 downto 23)) - ("00" & Y(30 downto 23));
   sR <= X(31) xor Y(31);
   -- early exception handling 
   exnXY <= X(33 downto 32) & Y(33 downto 32);
   with exnXY select
      exnR0 <= 
         "01"  when "0101",                   -- normal
         "00"  when "0001" | "0010" | "0110", -- zero
         "10"  when "0100" | "1000" | "1001", -- overflow
         "11"  when others;                   -- NaN
    -- Prescaling
   with partialFY (22 downto 21) select
      fY <= 
         ("0" & partialFY & "0") + (partialFY & "00") when "00",
         ("00" & partialFY) + (partialFY & "00") when "01",
         partialFY &"00" when others;
   with partialFY (22 downto 21) select
      fX <= 
         ("00" & partialFX & "0") + ("0" & partialFX & "00") when "00",
         ("000" & partialFX) + ("0" & partialFX & "00") when "01",
         "0" & partialFX &"00" when others;
   w9 <=  "00" & fX;
   ----------------Synchro barrier, entering cycle 1----------------
   sel9 <= w9_d1(28 downto 24) & fY_d1(23 downto 22);
   SelFunctionTable9: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel9,
                 Y => q9);
   w9pad <= w9_d1 & '0';
   with q9(1 downto 0) select 
   w8fulla <= 
      w9pad - ("0000" & fY_d1)			when "01",
      w9pad + ("0000" & fY_d1)			when "11",
      w9pad + ("000" & fY_d1 & "0")	  when "10",
      w9pad 			   		  when others;
   with q9(3 downto 1) select 
   fYdec8 <= 
      ("00" & fY_d1 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d1 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q9(3) select
   w8full <= 
      w8fulla - fYdec8			when '0',
      w8fulla + fYdec8			when others;
   w8 <= w8full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 2----------------
   sel8 <= w8_d1(28 downto 24) & fY_d2(23 downto 22);
   SelFunctionTable8: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel8,
                 Y => q8);
   w8pad <= w8_d1 & '0';
   with q8(1 downto 0) select 
   w7fulla <= 
      w8pad - ("0000" & fY_d2)			when "01",
      w8pad + ("0000" & fY_d2)			when "11",
      w8pad + ("000" & fY_d2 & "0")	  when "10",
      w8pad 			   		  when others;
   with q8(3 downto 1) select 
   fYdec7 <= 
      ("00" & fY_d2 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d2 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q8(3) select
   w7full <= 
      w7fulla - fYdec7			when '0',
      w7fulla + fYdec7			when others;
   w7 <= w7full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 3----------------
   sel7 <= w7_d1(28 downto 24) & fY_d3(23 downto 22);
   SelFunctionTable7: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel7,
                 Y => q7);
   w7pad <= w7_d1 & '0';
   with q7(1 downto 0) select 
   w6fulla <= 
      w7pad - ("0000" & fY_d3)			when "01",
      w7pad + ("0000" & fY_d3)			when "11",
      w7pad + ("000" & fY_d3 & "0")	  when "10",
      w7pad 			   		  when others;
   with q7(3 downto 1) select 
   fYdec6 <= 
      ("00" & fY_d3 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d3 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q7(3) select
   w6full <= 
      w6fulla - fYdec6			when '0',
      w6fulla + fYdec6			when others;
   w6 <= w6full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 4----------------
   sel6 <= w6_d1(28 downto 24) & fY_d4(23 downto 22);
   SelFunctionTable6: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel6,
                 Y => q6);
   w6pad <= w6_d1 & '0';
   with q6(1 downto 0) select 
   w5fulla <= 
      w6pad - ("0000" & fY_d4)			when "01",
      w6pad + ("0000" & fY_d4)			when "11",
      w6pad + ("000" & fY_d4 & "0")	  when "10",
      w6pad 			   		  when others;
   with q6(3 downto 1) select 
   fYdec5 <= 
      ("00" & fY_d4 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d4 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q6(3) select
   w5full <= 
      w5fulla - fYdec5			when '0',
      w5fulla + fYdec5			when others;
   w5 <= w5full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 5----------------
   sel5 <= w5_d1(28 downto 24) & fY_d5(23 downto 22);
   SelFunctionTable5: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel5,
                 Y => q5);
   w5pad <= w5_d1 & '0';
   with q5(1 downto 0) select 
   w4fulla <= 
      w5pad - ("0000" & fY_d5)			when "01",
      w5pad + ("0000" & fY_d5)			when "11",
      w5pad + ("000" & fY_d5 & "0")	  when "10",
      w5pad 			   		  when others;
   with q5(3 downto 1) select 
   fYdec4 <= 
      ("00" & fY_d5 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d5 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q5(3) select
   w4full <= 
      w4fulla - fYdec4			when '0',
      w4fulla + fYdec4			when others;
   w4 <= w4full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 6----------------
   sel4 <= w4_d1(28 downto 24) & fY_d6(23 downto 22);
   SelFunctionTable4: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel4,
                 Y => q4);
   w4pad <= w4_d1 & '0';
   with q4(1 downto 0) select 
   w3fulla <= 
      w4pad - ("0000" & fY_d6)			when "01",
      w4pad + ("0000" & fY_d6)			when "11",
      w4pad + ("000" & fY_d6 & "0")	  when "10",
      w4pad 			   		  when others;
   with q4(3 downto 1) select 
   fYdec3 <= 
      ("00" & fY_d6 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d6 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q4(3) select
   w3full <= 
      w3fulla - fYdec3			when '0',
      w3fulla + fYdec3			when others;
   w3 <= w3full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 7----------------
   sel3 <= w3_d1(28 downto 24) & fY_d7(23 downto 22);
   SelFunctionTable3: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel3,
                 Y => q3);
   w3pad <= w3_d1 & '0';
   with q3(1 downto 0) select 
   w2fulla <= 
      w3pad - ("0000" & fY_d7)			when "01",
      w3pad + ("0000" & fY_d7)			when "11",
      w3pad + ("000" & fY_d7 & "0")	  when "10",
      w3pad 			   		  when others;
   with q3(3 downto 1) select 
   fYdec2 <= 
      ("00" & fY_d7 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d7 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q3(3) select
   w2full <= 
      w2fulla - fYdec2			when '0',
      w2fulla + fYdec2			when others;
   w2 <= w2full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 8----------------
   sel2 <= w2_d1(28 downto 24) & fY_d8(23 downto 22);
   SelFunctionTable2: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel2,
                 Y => q2);
   w2pad <= w2_d1 & '0';
   with q2(1 downto 0) select 
   w1fulla <= 
      w2pad - ("0000" & fY_d8)			when "01",
      w2pad + ("0000" & fY_d8)			when "11",
      w2pad + ("000" & fY_d8 & "0")	  when "10",
      w2pad 			   		  when others;
   with q2(3 downto 1) select 
   fYdec1 <= 
      ("00" & fY_d8 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d8 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q2(3) select
   w1full <= 
      w1fulla - fYdec1			when '0',
      w1fulla + fYdec1			when others;
   w1 <= w1full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 9----------------
   sel1 <= w1_d1(28 downto 24) & fY_d9(23 downto 22);
   SelFunctionTable1: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel1,
                 Y => q1);
   w1pad <= w1_d1 & '0';
   with q1(1 downto 0) select 
   w0fulla <= 
      w1pad - ("0000" & fY_d9)			when "01",
      w1pad + ("0000" & fY_d9)			when "11",
      w1pad + ("000" & fY_d9 & "0")	  when "10",
      w1pad 			   		  when others;
   with q1(3 downto 1) select 
   fYdec0 <= 
      ("00" & fY_d9 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d9 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q1(3) select
   w0full <= 
      w0fulla - fYdec0			when '0',
      w0fulla + fYdec0			when others;
   w0 <= w0full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 10----------------
   q0(3 downto 0) <= "0000" when  w0_d1 = (28 downto 0 => '0')
                else w0_d1(28) & "010";
   qP9 <=      q9_d9(2 downto 0);
   qM9 <=      q9_d9(3) & "00";
   qP8 <=      q8_d8(2 downto 0);
   qM8 <=      q8_d8(3) & "00";
   qP7 <=      q7_d7(2 downto 0);
   qM7 <=      q7_d7(3) & "00";
   qP6 <=      q6_d6(2 downto 0);
   qM6 <=      q6_d6(3) & "00";
   qP5 <=      q5_d5(2 downto 0);
   qM5 <=      q5_d5(3) & "00";
   qP4 <=      q4_d4(2 downto 0);
   qM4 <=      q4_d4(3) & "00";
   qP3 <=      q3_d3(2 downto 0);
   qM3 <=      q3_d3(3) & "00";
   qP2 <=      q2_d2(2 downto 0);
   qM2 <=      q2_d2(3) & "00";
   qP1 <=      q1_d1(2 downto 0);
   qM1 <=      q1_d1(3) & "00";
   qP0 <= q0(2 downto 0);
   qM0 <= q0(3)  & "00";
   qP <= qP9 & qP8 & qP7 & qP6 & qP5 & qP4 & qP3 & qP2 & qP1 & qP0;
   qM <= qM9(1 downto 0) & qM8 & qM7 & qM6 & qM5 & qM4 & qM3 & qM2 & qM1 & qM0 & "0";
   fR0 <= qP - qM;
   ----------------Synchro barrier, entering cycle 11----------------
   fR <= fR0_d1(29 downto 2) & (fR0_d1(0) or fR0_d1(1)); 
   -- normalisation
   with fR(27) select
      fRn1 <= fR(27 downto 2) & (fR(0) or fR(1)) when '1',
              fR(26 downto 0)          when others;
   expR1 <= expR0_d11 + ("000" & (6 downto 1 => '1') & fR(27)); -- add back bias
   round <= fRn1(2) and (fRn1(0) or fRn1(1) or fRn1(3)); -- fRn1(0) is the sticky bit
   ----------------Synchro barrier, entering cycle 12----------------
   -- final rounding
   expfrac <= expR1_d1 & fRn1_d1(25 downto 3) ;
   expfracR <= expfrac + ((32 downto 1 => '0') & round_d1);
   exnR <=      "00"  when expfracR(32) = '1'   -- underflow
           else "10"  when  expfracR(32 downto 31) =  "01" -- overflow
           else "01";      -- 00, normal case
   with exnR0_d12 select
      exnRfinal <= 
         exnR   when "01", -- normal
         exnR0_d12  when others;
   R <= exnRfinal & sR_d12 & expfracR(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_348_mult_8en9_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_348_mult_8en9_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_348_mult_8en9_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100110110001110101101010011000001";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_125_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 125 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_125_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_125_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      Y <= s124;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 52 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      Y <= s51;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 47 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      Y <= s46;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 63 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      Y <= s62;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 37 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      Y <= s36;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_71_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 71 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_71_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_71_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      Y <= s70;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 68 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      Y <= s67;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 43 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      Y <= s42;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 23 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      Y <= s22;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 49 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      Y <= s48;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 55 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      Y <= s54;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 54 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      Y <= s53;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 35 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      Y <= s34;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 34 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      Y <= s33;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 41 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      Y <= s40;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 46 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      Y <= s45;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 53 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      Y <= s52;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      Y <= s15;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 24 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      Y <= s23;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 28 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      Y <= s27;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 22 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      Y <= s21;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 65 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      Y <= s64;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 48 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      Y <= s47;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 30 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      Y <= s29;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 31 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      Y <= s30;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 44 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      Y <= s43;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "001" when "0101",
      "000" when "0110",
      "000" when "0111",
      "010" when "1000",
      "000" when "1001",
      "000" when "1010",
      "011" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when "1110",
      "100" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when "1110",
      "000" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when "1110",
      "000" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when "1110",
      "000" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when "1110",
      "000" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when "1110",
      "000" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when "1110",
      "000" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "001" when "0101",
      "000" when "0110",
      "000" when "0111",
      "010" when "1000",
      "000" when "1001",
      "000" when "1010",
      "011" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when "1110",
      "100" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when "1110",
      "000" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "001" when "0010",
      "000" when "0011",
      "000" when "0100",
      "010" when "0101",
      "000" when "0110",
      "000" when "0111",
      "011" when "1000",
      "000" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when "1110",
      "100" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when "1110",
      "000" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when "1110",
      "000" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add17_4_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add17_4_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add17_4_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0001" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0100" when "0011",
      "0000" when "0100",
      "0111" when "0101",
      "0010" when "0110",
      "0000" when "0111",
      "1010" when "1000",
      "0101" when "1001",
      "0000" when "1010",
      "0110" when "1011",
      "0011" when "1100",
      "0000" when "1101",
      "1001" when "1110",
      "1000" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add17_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add17_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add17_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Add17_4_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add17_4_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add17_4_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add17_4_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add17_4_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0001" when "0000",
      "0000" when "0001",
      "1010" when "0010",
      "0111" when "0011",
      "0000" when "0100",
      "0000" when "0101",
      "0010" when "0110",
      "0000" when "0111",
      "0011" when "1000",
      "0101" when "1001",
      "0000" when "1010",
      "1000" when "1011",
      "0100" when "1100",
      "0000" when "1101",
      "1001" when "1110",
      "0110" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add17_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add17_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add17_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Add17_4_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add17_4_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add51_4_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add51_4_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add51_4_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0110" when "0000",
      "0000" when "0001",
      "0001" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0100" when "0101",
      "0010" when "0110",
      "0000" when "0111",
      "0011" when "1000",
      "1000" when "1001",
      "0000" when "1010",
      "0111" when "1011",
      "0000" when "1100",
      "0000" when "1101",
      "0101" when "1110",
      "1001" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add51_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add51_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add51_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Add51_4_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add51_4_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add51_4_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add51_4_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add51_4_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0101" when "0000",
      "0000" when "0001",
      "1001" when "0010",
      "1000" when "0011",
      "0000" when "0100",
      "0110" when "0101",
      "0000" when "0110",
      "0000" when "0111",
      "0010" when "1000",
      "0011" when "1001",
      "0000" when "1010",
      "0100" when "1011",
      "0000" when "1100",
      "0000" when "1101",
      "0111" when "1110",
      "0001" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add51_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add51_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add51_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Add51_4_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add51_4_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product105_4_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product105_4_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product105_4_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "1001" when "0001",
      "0101" when "0010",
      "0000" when "0011",
      "1010" when "0100",
      "0001" when "0101",
      "0000" when "0110",
      "0011" when "0111",
      "1000" when "1000",
      "0000" when "1001",
      "0111" when "1010",
      "0100" when "1011",
      "0010" when "1100",
      "0000" when "1101",
      "0000" when "1110",
      "0110" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product105_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product105_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product105_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product105_4_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product105_4_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product105_4_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product105_4_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product105_4_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "0111" when "0001",
      "0101" when "0010",
      "0000" when "0011",
      "1000" when "0100",
      "0010" when "0101",
      "0000" when "0110",
      "1001" when "0111",
      "0011" when "1000",
      "0000" when "1001",
      "0001" when "1010",
      "0100" when "1011",
      "0110" when "1100",
      "0000" when "1101",
      "0000" when "1110",
      "1010" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product105_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product105_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product105_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product105_4_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product105_4_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product512_4_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product512_4_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product512_4_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "1010" when "0001",
      "0111" when "0010",
      "0000" when "0011",
      "1001" when "0100",
      "0011" when "0101",
      "0000" when "0110",
      "1000" when "0111",
      "0000" when "1000",
      "0000" when "1001",
      "0110" when "1010",
      "0101" when "1011",
      "0100" when "1100",
      "0000" when "1101",
      "0010" when "1110",
      "0001" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product512_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product512_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product512_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product512_4_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product512_4_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product512_4_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product512_4_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product512_4_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "0101" when "0001",
      "1010" when "0010",
      "0000" when "0011",
      "0110" when "0100",
      "0000" when "0101",
      "0000" when "0110",
      "0001" when "0111",
      "0100" when "1000",
      "0000" when "1001",
      "1001" when "1010",
      "1000" when "1011",
      "0111" when "1100",
      "0000" when "1101",
      "0010" when "1110",
      "0011" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product512_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product512_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product512_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product512_4_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product512_4_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product55_4_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product55_4_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product55_4_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "1010" when "0001",
      "0110" when "0010",
      "0000" when "0011",
      "0011" when "0100",
      "0010" when "0101",
      "0000" when "0110",
      "1001" when "0111",
      "0111" when "1000",
      "0000" when "1001",
      "1000" when "1010",
      "0101" when "1011",
      "0100" when "1100",
      "0000" when "1101",
      "0000" when "1110",
      "0001" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product55_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product55_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product55_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product55_4_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product55_4_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product55_4_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product55_4_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product55_4_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "0111" when "0001",
      "1010" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0011" when "0101",
      "0000" when "0110",
      "0110" when "0111",
      "0101" when "1000",
      "0000" when "1001",
      "0100" when "1010",
      "1001" when "1011",
      "1000" when "1100",
      "0000" when "1101",
      "0010" when "1110",
      "0001" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product55_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product55_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product55_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product55_4_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product55_4_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product611_4_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product611_4_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product611_4_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "1010" when "0001",
      "1001" when "0010",
      "0000" when "0011",
      "0100" when "0100",
      "0011" when "0101",
      "0000" when "0110",
      "0111" when "0111",
      "0000" when "1000",
      "0000" when "1001",
      "1000" when "1010",
      "0110" when "1011",
      "0101" when "1100",
      "0000" when "1101",
      "0001" when "1110",
      "0010" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product611_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product611_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product611_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product611_4_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product611_4_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product611_4_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product611_4_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product611_4_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "0110" when "0001",
      "0101" when "0010",
      "0000" when "0011",
      "0111" when "0100",
      "0000" when "0101",
      "0000" when "0110",
      "1000" when "0111",
      "0001" when "1000",
      "0000" when "1001",
      "0010" when "1010",
      "1001" when "1011",
      "0100" when "1100",
      "0000" when "1101",
      "0011" when "1110",
      "1010" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product611_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product611_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product611_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product611_4_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product611_4_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "1000" when "0001",
      "0111" when "0010",
      "0000" when "0011",
      "0100" when "0100",
      "0011" when "0101",
      "0000" when "0110",
      "0000" when "0111",
      "0001" when "1000",
      "0000" when "1001",
      "0110" when "1010",
      "0101" when "1011",
      "0000" when "1100",
      "0000" when "1101",
      "0010" when "1110",
      "0000" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "0110" when "0001",
      "0101" when "0010",
      "0000" when "0011",
      "0111" when "0100",
      "0000" when "0101",
      "0000" when "0110",
      "0010" when "0111",
      "0001" when "1000",
      "0000" when "1001",
      "0011" when "1010",
      "0100" when "1011",
      "0000" when "1100",
      "0000" when "1101",
      "1000" when "1110",
      "0000" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Subtract12_3_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract12_3_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract12_3_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "0101" when "0001",
      "0100" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0110" when "0101",
      "0000" when "0110",
      "1010" when "0111",
      "0001" when "1000",
      "1011" when "1001",
      "0010" when "1010",
      "0111" when "1011",
      "1001" when "1100",
      "0000" when "1101",
      "0011" when "1110",
      "1000" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract12_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract12_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract12_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract12_3_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Subtract12_3_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Subtract12_3_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract12_3_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract12_3_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "1001" when "0001",
      "0001" when "0010",
      "0000" when "0011",
      "0110" when "0100",
      "1010" when "0101",
      "0000" when "0110",
      "0101" when "0111",
      "0111" when "1000",
      "1011" when "1001",
      "1000" when "1010",
      "0010" when "1011",
      "0100" when "1100",
      "0000" when "1101",
      "0000" when "1110",
      "0011" when "1111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract12_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract12_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract12_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract12_3_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Subtract12_3_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Subtract10_4_impl_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract10_4_impl_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract10_4_impl_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "010" when "0100",
      "000" when "0101",
      "000" when "0110",
      "100" when "0111",
      "000" when "1000",
      "000" when "1001",
      "000" when "1010",
      "011" when "1011",
      "000" when "1100",
      "000" when "1101",
      "001" when "1110",
      "000" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract10_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract10_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract10_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract10_4_impl_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Subtract10_4_impl_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Subtract10_4_impl_1_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract10_4_impl_1_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract10_4_impl_1_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "011" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "010" when "0111",
      "000" when "1000",
      "000" when "1001",
      "000" when "1010",
      "001" when "1011",
      "000" when "1100",
      "000" when "1101",
      "100" when "1110",
      "000" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract10_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract10_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract10_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract10_4_impl_1_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Subtract10_4_impl_1_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "001" when "0011",
      "000" when "0100",
      "000" when "0101",
      "010" when "0110",
      "000" when "0111",
      "000" when "1000",
      "011" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when "1100",
      "100" when "1101",
      "000" when "1110",
      "000" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "001" when "0011",
      "000" when "0100",
      "000" when "0101",
      "010" when "0110",
      "000" when "0111",
      "000" when "1000",
      "011" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when "1100",
      "100" when "1101",
      "000" when "1110",
      "000" when "1111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 99 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      Y <= s98;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_98_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 98 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_98_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_98_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      Y <= s97;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_123_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 123 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_123_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_123_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      Y <= s122;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_108_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 108 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_108_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_108_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      Y <= s107;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_94_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 94 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_94_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_94_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      Y <= s93;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_119_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 119 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_119_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_119_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      Y <= s118;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 104 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      Y <= s103;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 107 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      Y <= s106;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      Y <= s17;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 26 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      Y <= s25;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 32 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      Y <= s31;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 50 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      Y <= s49;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 27 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      Y <= s26;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 61 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      Y <= s60;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      Y <= s18;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 64 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      Y <= s63;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 62 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      Y <= s61;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_144_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 144 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_144_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_144_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      Y <= s143;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          Ldiff_UU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1_0 : in std_logic_vector(31 downto 0);
          R_U_0 : in std_logic_vector(31 downto 0);
          R_V_0 : in std_logic_vector(31 downto 0);
          R_W_0 : in std_logic_vector(31 downto 0);
          Inv_11_0 : out std_logic_vector(31 downto 0);
          Inv_12_0 : out std_logic_vector(31 downto 0);
          Inv_13_0 : out std_logic_vector(31 downto 0);
          Inv_21_0 : out std_logic_vector(31 downto 0);
          Inv_22_0 : out std_logic_vector(31 downto 0);
          Inv_23_0 : out std_logic_vector(31 downto 0);
          Inv_31_0 : out std_logic_vector(31 downto 0);
          Inv_32_0 : out std_logic_vector(31 downto 0);
          Inv_33_0 : out std_logic_vector(31 downto 0);
          Inv_41_0 : out std_logic_vector(31 downto 0);
          Inv_42_0 : out std_logic_vector(31 downto 0);
          Inv_43_0 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_16_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(3 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_16_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_5_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_11_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_10_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_9_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_12_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_348_mult_8en9_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_125_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_71_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add17_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add17_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add51_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add51_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product105_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product105_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product512_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product512_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product55_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product55_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product611_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product611_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract12_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract12_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract10_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract10_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_98_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_123_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_108_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_94_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_119_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_144_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount161_out : std_logic_vector(3 downto 0) := (others => '0');
signal Ldiff_UU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_11_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_12_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_13_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_21_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_22_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_23_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_31_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_32_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_33_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_41_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_42_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_43_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add101_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add141_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add151_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add151_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add151_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add151_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add151_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add151_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add16_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add17_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add17_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add17_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add24_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add24_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add24_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add51_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add51_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add51_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product112_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product112_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product112_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product113_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product102_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product102_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product102_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product104_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product104_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product104_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product104_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product104_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product104_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product104_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product104_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product104_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product105_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product105_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product105_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product105_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product105_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product105_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product105_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product105_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product105_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product241_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product241_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product241_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product361_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product361_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product361_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product391_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product391_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product391_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product441_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product441_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product441_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product491_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product491_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product491_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product512_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product56_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product56_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product56_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product611_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product611_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product611_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product611_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product611_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product611_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product811_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product811_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product811_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract10_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Divide_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Divide_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Divide_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay131No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay125No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay21No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay33No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay33No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay67No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay67No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay35No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay35No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay35No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_11_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_12_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_13_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_21_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_22_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_23_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_31_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_32_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_33_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_41_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_42_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_43_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Add17_4_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Add17_4_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Add51_4_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Add51_4_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product105_4_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product105_4_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product512_4_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product512_4_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product55_4_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product55_4_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product611_4_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product611_4_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product811_4_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product811_4_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Subtract12_3_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Subtract12_3_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Subtract10_4_impl_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Subtract10_4_impl_1_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Divide_0_impl_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Divide_0_impl_1_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out_to_Product108_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out_to_Product108_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out_to_Product108_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out_to_Product108_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out_to_Product110_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out_to_Product110_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out_to_Product109_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out_to_Product109_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out_to_Product109_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out_to_Product109_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No2_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out_to_Product111_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out_to_Product111_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out_to_Product210_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out_to_Product210_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out_to_Product210_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out_to_Product210_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No1_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No1_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out_to_Product210_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out_to_Product210_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No2_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out_to_Product210_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out_to_Product210_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No3_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out_to_Product210_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Product210_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No4_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No4_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No5_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No6_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No7_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Product310_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Product310_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Product310_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Product310_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay133No9_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Product610_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Product610_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No30_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No16_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Product610_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Product610_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Product610_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Product610_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Product610_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Product610_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay131No4_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Product810_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Product810_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Product810_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Product810_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Product810_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Product810_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay125No3_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Product810_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Product810_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_11_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_12_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_13_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_21_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_22_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_23_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_31_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_32_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_33_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_41_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_42_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_43_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Add30_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Add30_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No3_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Add30_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Add30_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No3_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No2_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Add110_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Add110_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No3_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay35No3_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Add101_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Add101_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No1_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No132_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Add121_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Add121_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No4_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No4_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Add141_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Add141_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No40_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay21No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No65_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Add151_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Add151_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay35No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No2_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Add151_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Add151_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No17_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay35No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No3_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay67No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Add16_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Add16_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay67No3_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No3_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No4_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No3_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Add17_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Add17_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No4_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No4_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No69_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Add24_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Add24_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No1_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Add51_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Add51_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No4_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No4_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No4_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Product112_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Product112_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Product112_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Product112_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Product112_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Product112_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Product113_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Product113_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Product102_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Product102_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No36_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Product102_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Product102_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Product102_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Product102_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No38_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Product104_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Product104_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Product104_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Product104_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Product104_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Product104_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Product105_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Product105_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Product105_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Product105_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Product105_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Product105_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Product241_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Product241_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Product321_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Product321_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Product361_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Product361_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Product391_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Product391_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Product441_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Product441_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Product491_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Product491_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Product512_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Product512_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Product55_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Product55_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out_to_Product56_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out_to_Product56_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out_to_Product611_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out_to_Product611_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out_to_Product611_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out_to_Product611_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No24_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out_to_Product811_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out_to_Product811_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay33No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay33No1_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No2_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No3_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out_to_Subtract12_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out_to_Subtract12_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No4_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out_to_Subtract10_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out_to_Subtract10_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No4_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount161_instance: ModuloCounter_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount161_out);
Ldiff_UU_del_1_0_IEEE <= Ldiff_UU_del_1_0;
   Ldiff_UU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_0_out,
                 X => Ldiff_UU_del_1_0_IEEE);
Ldiff_UV_del_1_0_IEEE <= Ldiff_UV_del_1_0;
   Ldiff_UV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_0_out,
                 X => Ldiff_UV_del_1_0_IEEE);
Ldiff_UW_del_1_0_IEEE <= Ldiff_UW_del_1_0;
   Ldiff_UW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_0_out,
                 X => Ldiff_UW_del_1_0_IEEE);
Ldiff_VU_del_1_0_IEEE <= Ldiff_VU_del_1_0;
   Ldiff_VU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_0_out,
                 X => Ldiff_VU_del_1_0_IEEE);
Ldiff_VV_del_1_0_IEEE <= Ldiff_VV_del_1_0;
   Ldiff_VV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_0_out,
                 X => Ldiff_VV_del_1_0_IEEE);
Ldiff_VW_del_1_0_IEEE <= Ldiff_VW_del_1_0;
   Ldiff_VW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_0_out,
                 X => Ldiff_VW_del_1_0_IEEE);
Ldiff_WU_del_1_0_IEEE <= Ldiff_WU_del_1_0;
   Ldiff_WU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_0_out,
                 X => Ldiff_WU_del_1_0_IEEE);
Ldiff_WV_del_1_0_IEEE <= Ldiff_WV_del_1_0;
   Ldiff_WV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_0_out,
                 X => Ldiff_WV_del_1_0_IEEE);
Ldiff_WW_del_1_0_IEEE <= Ldiff_WW_del_1_0;
   Ldiff_WW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_0_out,
                 X => Ldiff_WW_del_1_0_IEEE);
R_U_0_IEEE <= R_U_0;
   R_U_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_0_out,
                 X => R_U_0_IEEE);
R_V_0_IEEE <= R_V_0;
   R_V_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_0_out,
                 X => R_V_0_IEEE);
R_W_0_IEEE <= R_W_0;
   R_W_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_0_out,
                 X => R_W_0_IEEE);

Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast <= Delay1No_out;
Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast <= Delay1No1_out;
   Product108_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_0_impl_out,
                 X => Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg1_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg560_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg175_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg175_out;
SharedReg564_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg89_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg89_out;
SharedReg42_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg42_out;
SharedReg143_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg143_out;
SharedReg40_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg40_out;
SharedReg93_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg93_out;
SharedReg220_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg220_out;
SharedReg556_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg557_out;
   MUX_Product108_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg143_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg40_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg93_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg220_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg556_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg557_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg175_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg89_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg42_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product108_0_impl_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_0_impl_0_out,
                 Y => Delay1No_out);

SharedReg254_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg254_out;
SharedReg20_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg560_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg10_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg10_out;
SharedReg22_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg22_out;
SharedReg367_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg367_out;
SharedReg34_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg34_out;
SharedReg369_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg369_out;
SharedReg576_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg576_out;
SharedReg257_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg257_out;
SharedReg257_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg257_out;
   MUX_Product108_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg254_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg367_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg34_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg369_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg576_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg257_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg257_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg10_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg22_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product108_0_impl_1_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_0_impl_1_out,
                 Y => Delay1No1_out);

Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast <= Delay1No2_out;
Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast <= Delay1No3_out;
   Product108_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_1_impl_out,
                 X => Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast);

SharedReg312_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg312_out;
SharedReg556_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg1_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg560_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg48_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg48_out;
SharedReg564_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg565_out;
SharedReg118_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg118_out;
SharedReg96_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg96_out;
SharedReg377_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg377_out;
SharedReg48_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg48_out;
SharedReg380_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg380_out;
   MUX_Product108_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg312_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg556_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg118_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg96_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg377_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg48_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg380_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg48_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product108_1_impl_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_1_impl_0_out,
                 Y => Delay1No2_out);

SharedReg24_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg24_out;
SharedReg266_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg266_out;
SharedReg266_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg266_out;
SharedReg264_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg264_out;
SharedReg20_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg560_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg565_out;
SharedReg16_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg16_out;
SharedReg11_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg11_out;
SharedReg23_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg23_out;
SharedReg5_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg5_out;
SharedReg337_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg337_out;
   MUX_Product108_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg24_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg266_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg16_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg11_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg23_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg5_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg337_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg266_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg264_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product108_1_impl_1_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_1_impl_1_out,
                 Y => Delay1No3_out);

Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast <= Delay1No4_out;
Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast <= Delay1No5_out;
   Product108_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_2_impl_out,
                 X => Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast);

SharedReg419_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg419_out;
SharedReg76_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg76_out;
SharedReg387_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg387_out;
SharedReg294_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg294_out;
SharedReg556_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg7_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg7_out;
SharedReg14_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg14_out;
SharedReg561_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg54_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg54_out;
SharedReg564_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg565_out;
SharedReg54_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg54_out;
SharedReg192_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg192_out;
   MUX_Product108_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg419_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg76_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg54_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg564_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg565_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg54_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg192_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg387_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg294_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg556_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg7_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg14_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product108_2_impl_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_2_impl_0_out,
                 Y => Delay1No4_out);

SharedReg567_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg5_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg345_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg345_out;
SharedReg24_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg24_out;
SharedReg298_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg298_out;
SharedReg298_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg298_out;
SharedReg351_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg351_out;
SharedReg13_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg561_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg565_out;
SharedReg32_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg22_out;
   MUX_Product108_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg564_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg565_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg32_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg22_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg345_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg24_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg298_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg298_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg351_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg13_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product108_2_impl_1_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_2_impl_1_out,
                 Y => Delay1No5_out);

Delay1No6_out_to_Product108_3_impl_parent_implementedSystem_port_0_cast <= Delay1No6_out;
Delay1No7_out_to_Product108_3_impl_parent_implementedSystem_port_1_cast <= Delay1No7_out;
   Product108_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_3_impl_out,
                 X => Delay1No6_out_to_Product108_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No7_out_to_Product108_3_impl_parent_implementedSystem_port_1_cast);

SharedReg565_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg106_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg106_out;
SharedReg61_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg61_out;
SharedReg471_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg471_out;
SharedReg231_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg231_out;
SharedReg85_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg85_out;
SharedReg286_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg286_out;
SharedReg556_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg7_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg7_out;
SharedReg14_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg14_out;
SharedReg561_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg60_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg60_out;
SharedReg564_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg564_out;
   MUX_Product108_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg106_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg7_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg14_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg60_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg564_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg61_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg471_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg231_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg85_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg286_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg556_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product108_3_impl_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_3_impl_0_out,
                 Y => Delay1No6_out);

SharedReg565_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg16_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg11_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg11_out;
SharedReg299_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg299_out;
SharedReg34_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg34_out;
SharedReg301_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg301_out;
SharedReg24_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg24_out;
SharedReg288_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg288_out;
SharedReg352_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg352_out;
SharedReg307_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg307_out;
SharedReg13_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg31_out;
SharedReg561_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg564_out;
   MUX_Product108_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg13_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg31_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg564_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg11_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg299_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg34_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg301_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg24_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg288_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg352_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg307_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product108_3_impl_1_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_3_impl_1_out,
                 Y => Delay1No7_out);

Delay1No8_out_to_Product108_4_impl_parent_implementedSystem_port_0_cast <= Delay1No8_out;
Delay1No9_out_to_Product108_4_impl_parent_implementedSystem_port_1_cast <= Delay1No9_out;
   Product108_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_4_impl_out,
                 X => Delay1No8_out_to_Product108_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No9_out_to_Product108_4_impl_parent_implementedSystem_port_1_cast);

SharedReg561_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg70_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg70_out;
SharedReg137_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg137_out;
SharedReg565_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg565_out;
SharedReg64_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg64_out;
SharedReg513_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg513_out;
SharedReg171_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg171_out;
SharedReg64_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg64_out;
SharedReg211_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg211_out;
SharedReg446_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg446_out;
SharedReg556_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg558_out;
SharedReg7_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg7_out;
SharedReg8_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg8_out;
   MUX_Product108_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg446_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg556_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg557_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg558_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg7_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg8_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg70_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg137_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg565_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg64_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg513_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg171_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg64_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg211_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product108_4_impl_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_4_impl_0_out,
                 Y => Delay1No8_out);

SharedReg561_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg565_out;
SharedReg10_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg10_out;
SharedReg566_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg566_out;
SharedReg372_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg372_out;
SharedReg34_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg34_out;
SharedReg361_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg361_out;
SharedReg576_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg576_out;
SharedReg308_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg308_out;
SharedReg323_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg323_out;
SharedReg358_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg358_out;
SharedReg13_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg13_out;
SharedReg26_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg26_out;
   MUX_Product108_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg576_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg308_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg323_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg358_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg13_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg26_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg563_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg565_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg10_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg566_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg372_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg34_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg361_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product108_4_impl_1_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_4_impl_1_out,
                 Y => Delay1No9_out);

Delay1No10_out_to_Product110_4_impl_parent_implementedSystem_port_0_cast <= Delay1No10_out;
Delay1No11_out_to_Product110_4_impl_parent_implementedSystem_port_1_cast <= Delay1No11_out;
   Product110_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_4_impl_out,
                 X => Delay1No10_out_to_Product110_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No11_out_to_Product110_4_impl_parent_implementedSystem_port_1_cast);

SharedReg561_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg209_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg209_out;
SharedReg64_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg64_out;
SharedReg28_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg28_out;
SharedReg301_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg301_out;
SharedReg139_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg139_out;
SharedReg479_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg479_out;
SharedReg70_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg70_out;
SharedReg210_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg210_out;
SharedReg39_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg39_out;
SharedReg38_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg38_out;
SharedReg557_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg558_out;
SharedReg1_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1_out;
SharedReg14_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg14_out;
   MUX_Product110_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg39_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg38_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg557_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg558_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg14_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg209_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg64_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg28_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg301_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg139_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg479_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg70_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg210_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product110_4_impl_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_4_impl_0_out,
                 Y => Delay1No10_out);

SharedReg561_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg299_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg299_out;
SharedReg300_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg300_out;
SharedReg575_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg575_out;
SharedReg578_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg578_out;
SharedReg570_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg570_out;
SharedReg373_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg373_out;
SharedReg559_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg325_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg325_out;
SharedReg322_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg322_out;
SharedReg20_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg20_out;
SharedReg31_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg31_out;
   MUX_Product110_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg325_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg322_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg20_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg31_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg563_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg299_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg300_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg575_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg578_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg570_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg373_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product110_4_impl_1_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_4_impl_1_out,
                 Y => Delay1No11_out);

Delay1No12_out_to_Product109_2_impl_parent_implementedSystem_port_0_cast <= Delay1No12_out;
Delay1No13_out_to_Product109_2_impl_parent_implementedSystem_port_1_cast <= Delay1No13_out;
   Product109_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_2_impl_out,
                 X => Delay1No12_out_to_Product109_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No13_out_to_Product109_2_impl_parent_implementedSystem_port_1_cast);

SharedReg483_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg483_out;
SharedReg385_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg385_out;
SharedReg79_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg79_out;
SharedReg504_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg504_out;
SharedReg39_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg39_out;
SharedReg38_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg38_out;
SharedReg558_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg1_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg560_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg76_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg76_out;
SharedReg564_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg565_out;
SharedReg100_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg100_out;
SharedReg55_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg55_out;
   MUX_Product109_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg483_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg385_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg76_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg564_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg565_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg100_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg55_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg79_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg504_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg39_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg38_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product109_2_impl_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_2_impl_0_out,
                 Y => Delay1No12_out);

SharedReg344_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg344_out;
SharedReg34_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg34_out;
SharedReg346_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg346_out;
SharedReg576_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg576_out;
SharedReg559_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg272_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg272_out;
SharedReg20_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg20_out;
SharedReg560_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg565_out;
SharedReg16_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg16_out;
SharedReg11_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg11_out;
   MUX_Product109_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg344_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg34_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg564_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg565_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg16_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg11_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg346_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg576_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg272_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg20_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product109_2_impl_1_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_2_impl_1_out,
                 Y => Delay1No13_out);

Delay1No14_out_to_Product109_3_impl_parent_implementedSystem_port_0_cast <= Delay1No14_out;
Delay1No15_out_to_Product109_3_impl_parent_implementedSystem_port_1_cast <= Delay1No15_out;
   Product109_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_3_impl_out,
                 X => Delay1No14_out_to_Product109_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No15_out_to_Product109_3_impl_parent_implementedSystem_port_1_cast);

SharedReg565_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg82_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg82_out;
SharedReg394_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg394_out;
SharedReg60_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg60_out;
SharedReg397_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg397_out;
SharedReg392_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg392_out;
SharedReg485_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg485_out;
SharedReg39_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg39_out;
SharedReg38_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg38_out;
SharedReg558_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg1_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg560_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg82_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg82_out;
SharedReg564_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg564_out;
   MUX_Product109_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg82_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg82_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg564_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg394_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg397_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg392_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg485_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg39_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg38_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product109_3_impl_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_3_impl_0_out,
                 Y => Delay1No14_out);

SharedReg565_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg10_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg10_out;
SharedReg22_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg22_out;
SharedReg33_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg33_out;
SharedReg578_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg578_out;
SharedReg570_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg570_out;
SharedReg576_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg576_out;
SharedReg559_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg281_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg281_out;
SharedReg20_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg560_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg564_out;
   MUX_Product109_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg564_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg22_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg33_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg578_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg570_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg576_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg281_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product109_3_impl_1_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_3_impl_1_out,
                 Y => Delay1No15_out);

Delay1No16_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast <= Delay1No16_out;
Delay1No17_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast <= Delay1No17_out;
   Product111_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_0_impl_out,
                 X => Delay1No16_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No17_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg7_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg7_out;
SharedReg14_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg14_out;
SharedReg561_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg40_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg40_out;
SharedReg564_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg142_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg142_out;
SharedReg114_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg114_out;
SharedReg40_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg40_out;
SharedReg89_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg89_out;
SharedReg44_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg44_out;
SharedReg329_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg329_out;
SharedReg556_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg557_out;
   MUX_Product111_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg40_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg89_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg44_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg329_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg556_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg557_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg14_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg40_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg142_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg114_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product111_0_impl_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_0_impl_0_out,
                 Y => Delay1No16_out);

SharedReg335_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg335_out;
SharedReg13_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg31_out;
SharedReg561_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg16_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg16_out;
SharedReg11_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg11_out;
SharedReg23_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg23_out;
SharedReg5_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg5_out;
SharedReg368_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg368_out;
SharedReg35_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg35_out;
SharedReg256_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg256_out;
SharedReg255_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg255_out;
   MUX_Product111_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg335_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg23_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg5_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg368_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg35_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg256_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg255_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg31_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg16_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg11_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product111_0_impl_1_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_0_impl_1_out,
                 Y => Delay1No17_out);

Delay1No18_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast <= Delay1No18_out;
Delay1No19_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast <= Delay1No19_out;
   Product111_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_1_impl_out,
                 X => Delay1No18_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No19_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast);

SharedReg312_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg312_out;
SharedReg556_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg7_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg7_out;
SharedReg14_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg14_out;
SharedReg561_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg95_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg95_out;
SharedReg564_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg565_out;
SharedReg95_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg95_out;
SharedReg224_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg224_out;
SharedReg224_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg224_out;
SharedReg95_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg95_out;
SharedReg186_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg186_out;
   MUX_Product111_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg312_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg556_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg95_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg224_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg224_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg95_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg186_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg7_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg14_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg95_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product111_1_impl_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_1_impl_0_out,
                 Y => Delay1No18_out);

SharedReg24_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg24_out;
SharedReg317_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg317_out;
SharedReg265_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg265_out;
SharedReg343_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg343_out;
SharedReg13_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg31_out;
SharedReg561_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg565_out;
SharedReg32_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg22_out;
SharedReg336_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg336_out;
SharedReg28_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg28_out;
SharedReg311_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg311_out;
   MUX_Product111_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg24_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg317_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg32_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg22_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg336_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg28_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg311_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg265_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg343_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg13_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg31_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product111_1_impl_1_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_1_impl_1_out,
                 Y => Delay1No19_out);

Delay1No20_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast <= Delay1No20_out;
Delay1No21_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast <= Delay1No21_out;
   Product111_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_2_impl_out,
                 X => Delay1No20_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No21_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast);

SharedReg344_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg344_out;
SharedReg54_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg54_out;
SharedReg158_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg158_out;
SharedReg294_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg294_out;
SharedReg556_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg20_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg20_out;
SharedReg8_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg54_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg54_out;
SharedReg77_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg77_out;
SharedReg123_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg123_out;
SharedReg99_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg99_out;
   MUX_Product111_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg344_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg54_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg54_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg77_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg123_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg99_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg158_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg294_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg556_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg20_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg8_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product111_2_impl_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_2_impl_0_out,
                 Y => Delay1No20_out);

SharedReg17_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg17_out;
SharedReg28_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg28_out;
SharedReg293_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg293_out;
SharedReg24_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg24_out;
SharedReg341_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg341_out;
SharedReg273_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg273_out;
Delay133No2_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_7_cast <= Delay133No2_out;
SharedReg30_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg30_out;
SharedReg26_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg564_out;
SharedReg9_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg9_out;
SharedReg21_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg21_out;
SharedReg11_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg11_out;
   MUX_Product111_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg17_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg28_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg564_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg9_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg21_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg11_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg293_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg24_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg341_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg273_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay133No2_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg30_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg26_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product111_2_impl_1_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_2_impl_1_out,
                 Y => Delay1No21_out);

Delay1No22_out_to_Product111_3_impl_parent_implementedSystem_port_0_cast <= Delay1No22_out;
Delay1No23_out_to_Product111_3_impl_parent_implementedSystem_port_1_cast <= Delay1No23_out;
   Product111_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_3_impl_out,
                 X => Delay1No22_out_to_Product111_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No23_out_to_Product111_3_impl_parent_implementedSystem_port_1_cast);

SharedReg565_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg60_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg60_out;
SharedReg201_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg201_out;
SharedReg400_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg400_out;
SharedReg419_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg419_out;
SharedReg395_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg395_out;
SharedReg286_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg286_out;
SharedReg556_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg20_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg8_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg60_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg60_out;
   MUX_Product111_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg60_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg8_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg60_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg201_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg400_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg419_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg395_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg286_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg556_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product111_3_impl_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_3_impl_0_out,
                 Y => Delay1No22_out);

SharedReg565_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg32_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg22_out;
SharedReg567_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg567_out;
SharedReg5_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg5_out;
SharedReg300_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg300_out;
SharedReg24_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg24_out;
SharedReg350_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg350_out;
SharedReg282_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg282_out;
SharedReg290_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg290_out;
SharedReg30_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg30_out;
SharedReg26_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg564_out;
   MUX_Product111_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg32_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg30_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg26_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg564_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg22_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg567_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg5_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg300_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg24_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg350_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg282_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg290_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product111_3_impl_1_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_3_impl_1_out,
                 Y => Delay1No23_out);

Delay1No24_out_to_Product210_0_impl_parent_implementedSystem_port_0_cast <= Delay1No24_out;
Delay1No25_out_to_Product210_0_impl_parent_implementedSystem_port_1_cast <= Delay1No25_out;
   Product210_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_0_impl_out,
                 X => Delay1No24_out_to_Product210_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No25_out_to_Product210_0_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg20_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg8_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg89_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg89_out;
SharedReg564_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg113_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg113_out;
SharedReg426_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg426_out;
SharedReg426_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg426_out;
SharedReg113_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg113_out;
SharedReg218_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg218_out;
SharedReg6_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg6_out;
SharedReg556_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg557_out;
   MUX_Product210_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg426_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg113_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg218_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg6_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg556_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg557_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg8_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg89_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg113_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg426_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product210_0_impl_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_0_impl_0_out,
                 Y => Delay1No24_out);

Delay133No_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_1_cast <= Delay133No_out;
SharedReg30_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg30_out;
SharedReg26_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg32_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg22_out;
SharedReg367_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg367_out;
SharedReg28_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg28_out;
SharedReg328_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg328_out;
SharedReg370_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg370_out;
SharedReg333_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg333_out;
Delay130No_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_16_cast <= Delay130No_out;
   MUX_Product210_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay133No_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg367_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg28_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg328_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg370_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg333_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay130No_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg26_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg32_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg22_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product210_0_impl_1_out);

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_0_impl_1_out,
                 Y => Delay1No25_out);

Delay1No26_out_to_Product210_1_impl_parent_implementedSystem_port_0_cast <= Delay1No26_out;
Delay1No27_out_to_Product210_1_impl_parent_implementedSystem_port_1_cast <= Delay1No27_out;
   Product210_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_1_impl_out,
                 X => Delay1No26_out_to_Product210_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No27_out_to_Product210_1_impl_parent_implementedSystem_port_1_cast);

SharedReg227_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg227_out;
SharedReg556_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg20_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg8_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg563_out;
SharedReg95_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg95_out;
SharedReg49_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg49_out;
SharedReg148_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg148_out;
SharedReg117_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg117_out;
SharedReg435_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg435_out;
SharedReg183_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg183_out;
SharedReg50_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg50_out;
   MUX_Product210_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg227_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg556_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg49_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg148_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg117_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg435_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg183_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg50_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg8_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg95_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product210_1_impl_0_out);

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_1_impl_0_out,
                 Y => Delay1No26_out);

SharedReg576_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg576_out;
SharedReg316_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg316_out;
Delay130No1_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_3_cast <= Delay130No1_out;
Delay133No1_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_4_cast <= Delay133No1_out;
SharedReg30_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg30_out;
SharedReg26_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg9_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg9_out;
SharedReg21_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg21_out;
SharedReg11_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg11_out;
SharedReg309_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg309_out;
SharedReg5_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg5_out;
SharedReg337_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg337_out;
   MUX_Product210_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg576_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg316_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg9_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg21_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg11_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg309_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg5_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg337_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => Delay130No1_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay133No1_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg30_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg26_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product210_1_impl_1_out);

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_1_impl_1_out,
                 Y => Delay1No27_out);

Delay1No28_out_to_Product210_2_impl_parent_implementedSystem_port_0_cast <= Delay1No28_out;
Delay1No29_out_to_Product210_2_impl_parent_implementedSystem_port_1_cast <= Delay1No29_out;
   Product210_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_2_impl_out,
                 X => Delay1No28_out_to_Product210_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No29_out_to_Product210_2_impl_parent_implementedSystem_port_1_cast);

SharedReg291_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg291_out;
SharedReg156_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg156_out;
SharedReg78_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg78_out;
SharedReg194_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg194_out;
SharedReg556_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg419_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg419_out;
SharedReg20_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg20_out;
SharedReg2_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg2_out;
SharedReg561_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg99_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg99_out;
SharedReg565_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg565_out;
SharedReg156_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg156_out;
SharedReg495_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg495_out;
   MUX_Product210_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg291_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg156_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg99_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg565_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg156_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg495_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg78_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg194_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg556_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg419_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg20_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg2_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product210_2_impl_0_out);

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_2_impl_0_out,
                 Y => Delay1No28_out);

SharedReg344_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg344_out;
SharedReg5_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg345_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg345_out;
SharedReg576_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg576_out;
SharedReg297_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg297_out;
Delay130No2_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_6_cast <= Delay130No2_out;
SharedReg571_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg571_out;
SharedReg25_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg25_out;
SharedReg26_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg565_out;
SharedReg27_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg27_out;
SharedReg575_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg575_out;
   MUX_Product210_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg344_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg564_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg565_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg27_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg575_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg345_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg576_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg297_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay130No2_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg571_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg25_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg26_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product210_2_impl_1_out);

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_2_impl_1_out,
                 Y => Delay1No29_out);

Delay1No30_out_to_Product210_3_impl_parent_implementedSystem_port_0_cast <= Delay1No30_out;
Delay1No31_out_to_Product210_3_impl_parent_implementedSystem_port_1_cast <= Delay1No31_out;
   Product210_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_3_impl_out,
                 X => Delay1No30_out_to_Product210_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No31_out_to_Product210_3_impl_parent_implementedSystem_port_1_cast);

SharedReg469_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg469_out;
SharedReg130_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
SharedReg105_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg105_out;
SharedReg299_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg299_out;
SharedReg449_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg449_out;
SharedReg164_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg164_out;
SharedReg203_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg203_out;
SharedReg556_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg458_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg458_out;
SharedReg20_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg2_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg2_out;
SharedReg561_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg105_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg105_out;
   MUX_Product210_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg469_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg2_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg105_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg105_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg299_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg449_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg164_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg203_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg556_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg458_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product210_3_impl_0_out);

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_3_impl_0_out,
                 Y => Delay1No30_out);

SharedReg15_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg15_out;
SharedReg21_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg21_out;
SharedReg11_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg11_out;
SharedReg17_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg17_out;
SharedReg28_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg28_out;
SharedReg285_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg285_out;
SharedReg576_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg576_out;
SharedReg306_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg306_out;
Delay130No3_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_9_cast <= Delay130No3_out;
SharedReg571_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg571_out;
SharedReg25_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg25_out;
SharedReg26_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg564_out;
   MUX_Product210_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg15_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg21_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg25_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg26_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg564_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg11_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg17_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg28_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg285_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg576_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg306_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay130No3_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg571_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product210_3_impl_1_out);

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_3_impl_1_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Product210_4_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Product210_4_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Product210_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_4_impl_out,
                 X => Delay1No32_out_to_Product210_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Product210_4_impl_parent_implementedSystem_port_1_cast);

SharedReg561_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg64_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg64_out;
SharedReg169_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg169_out;
SharedReg565_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg565_out;
SharedReg470_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg470_out;
SharedReg464_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg464_out;
SharedReg400_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg400_out;
SharedReg137_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg137_out;
SharedReg244_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg244_out;
SharedReg362_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg362_out;
SharedReg556_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg558_out;
SharedReg20_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg20_out;
SharedReg2_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg2_out;
   MUX_Product210_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg362_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg556_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg557_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg558_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg20_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg2_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg64_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg169_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg565_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg470_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg464_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg400_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg137_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg244_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product210_4_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_4_impl_0_out,
                 Y => Delay1No32_out);

SharedReg561_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg565_out;
SharedReg16_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg16_out;
SharedReg566_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg566_out;
SharedReg23_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg23_out;
SharedReg5_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg5_out;
SharedReg29_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg29_out;
SharedReg35_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg35_out;
SharedReg324_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg324_out;
Delay130No4_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_13_cast <= Delay130No4_out;
Delay133No4_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_14_cast <= Delay133No4_out;
SharedReg30_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg30_out;
SharedReg26_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg26_out;
   MUX_Product210_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg35_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg324_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay130No4_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay133No4_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg30_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg26_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg563_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg565_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg16_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg566_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg23_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg5_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg29_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product210_4_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_4_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Product310_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_0_impl_out,
                 X => Delay1No34_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast);

SharedReg407_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg407_out;
SharedReg20_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg2_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg561_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg89_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg89_out;
SharedReg41_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg41_out;
SharedReg175_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg175_out;
SharedReg141_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg141_out;
SharedReg409_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg409_out;
SharedReg215_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg215_out;
SharedReg91_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg91_out;
SharedReg329_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg329_out;
SharedReg145_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg145_out;
SharedReg557_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg557_out;
   MUX_Product310_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg407_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg409_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg215_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg91_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg329_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg145_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg557_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg2_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg89_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg41_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg175_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg141_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product310_0_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_0_impl_0_out,
                 Y => Delay1No34_out);

SharedReg571_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg571_out;
SharedReg25_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg25_out;
SharedReg26_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg9_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg9_out;
SharedReg21_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg21_out;
SharedReg11_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg11_out;
SharedReg326_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg326_out;
SharedReg5_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg5_out;
SharedReg368_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg368_out;
SharedReg370_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg370_out;
SharedReg577_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg577_out;
Delay133No5_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_16_cast <= Delay133No5_out;
   MUX_Product310_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg571_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg25_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg326_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg5_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg368_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg370_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg577_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay133No5_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg26_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg9_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg21_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg11_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product310_0_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_0_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Product310_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_1_impl_out,
                 X => Delay1No36_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast);

SharedReg312_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg312_out;
SharedReg530_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg530_out;
SharedReg557_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg433_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg433_out;
SharedReg20_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg2_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg2_out;
SharedReg561_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg563_out;
SharedReg117_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg117_out;
SharedReg565_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg565_out;
SharedReg183_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg183_out;
SharedReg509_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg509_out;
SharedReg95_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg95_out;
SharedReg223_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg223_out;
SharedReg150_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg150_out;
   MUX_Product310_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg312_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg530_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg183_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg509_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg95_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg223_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg150_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg433_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg2_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg117_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product310_1_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_1_impl_0_out,
                 Y => Delay1No36_out);

SharedReg35_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg35_out;
SharedReg577_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg577_out;
Delay133No6_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast <= Delay133No6_out;
SharedReg571_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg571_out;
SharedReg25_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg25_out;
SharedReg26_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg565_out;
SharedReg27_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg27_out;
SharedReg575_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg575_out;
SharedReg33_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg33_out;
SharedReg310_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg310_out;
SharedReg337_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg337_out;
   MUX_Product310_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg35_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg577_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg27_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg575_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg33_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg310_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg337_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => Delay133No6_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg571_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg25_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg26_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product310_1_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_1_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Product310_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_2_impl_out,
                 X => Delay1No38_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast);

SharedReg231_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg231_out;
SharedReg191_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg191_out;
SharedReg125_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg125_out;
SharedReg294_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg294_out;
SharedReg389_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg389_out;
SharedReg557_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg449_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg449_out;
SharedReg1_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg99_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg99_out;
SharedReg123_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg123_out;
SharedReg565_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg565_out;
SharedReg232_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg232_out;
SharedReg419_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg419_out;
   MUX_Product310_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg231_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg191_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg99_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg123_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg565_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg232_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg419_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg125_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg294_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg389_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg449_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg8_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product310_2_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_2_impl_0_out,
                 Y => Delay1No38_out);

SharedReg567_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg292_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg292_out;
SharedReg345_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg345_out;
SharedReg35_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg35_out;
SharedReg577_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg577_out;
Delay133No7_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_6_cast <= Delay133No7_out;
SharedReg571_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg571_out;
SharedReg13_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg561_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg565_out;
SharedReg16_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg16_out;
SharedReg566_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg566_out;
   MUX_Product310_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg292_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg564_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg565_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg16_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg566_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg345_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg35_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg577_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay133No7_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg571_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg13_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product310_2_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_2_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Product310_3_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Product310_3_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Product310_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_3_impl_out,
                 X => Delay1No40_out_to_Product310_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Product310_3_impl_parent_implementedSystem_port_1_cast);

SharedReg239_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg239_out;
SharedReg163_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg163_out;
SharedReg454_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg454_out;
SharedReg283_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg283_out;
SharedReg82_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg82_out;
SharedReg84_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg84_out;
SharedReg286_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg286_out;
SharedReg398_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg398_out;
SharedReg557_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg469_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg469_out;
SharedReg1_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg105_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg105_out;
SharedReg130_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg130_out;
   MUX_Product310_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg239_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg163_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg8_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg105_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg130_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg454_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg283_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg82_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg84_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg286_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg398_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg469_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product310_3_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_3_impl_0_out,
                 Y => Delay1No40_out);

SharedReg574_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg574_out;
SharedReg27_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg27_out;
SharedReg575_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg575_out;
SharedReg299_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg299_out;
SharedReg5_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg5_out;
SharedReg300_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg300_out;
SharedReg35_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg35_out;
SharedReg577_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg577_out;
SharedReg290_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg290_out;
SharedReg571_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg571_out;
SharedReg13_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg31_out;
SharedReg561_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg564_out;
   MUX_Product310_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg574_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg13_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg31_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg564_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg575_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg299_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg5_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg300_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg35_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg577_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg290_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg571_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product310_3_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_3_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Product310_4_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Product310_4_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Product310_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_4_impl_out,
                 X => Delay1No42_out_to_Product310_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Product310_4_impl_parent_implementedSystem_port_1_cast);

SharedReg561_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg563_out;
SharedReg209_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg209_out;
SharedReg565_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg565_out;
SharedReg137_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg137_out;
SharedReg516_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg516_out;
SharedReg441_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg441_out;
SharedReg169_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg169_out;
SharedReg18_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg18_out;
SharedReg6_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg6_out;
SharedReg556_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg557_out;
SharedReg169_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg169_out;
SharedReg20_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg20_out;
SharedReg8_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg8_out;
   MUX_Product310_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg6_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg556_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg557_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg169_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg20_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg8_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg563_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg209_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg565_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg137_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg516_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg441_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg169_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg18_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product310_4_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_4_impl_0_out,
                 Y => Delay1No42_out);

SharedReg561_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg565_out;
SharedReg32_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg32_out;
SharedReg566_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg566_out;
SharedReg372_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg372_out;
SharedReg28_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg28_out;
SharedReg374_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg374_out;
SharedReg375_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg375_out;
SharedReg365_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg365_out;
Delay133No9_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_13_cast <= Delay133No9_out;
SharedReg571_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg571_out;
SharedReg25_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg25_out;
SharedReg31_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg31_out;
   MUX_Product310_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg375_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg365_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay133No9_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg571_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg25_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg31_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg563_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg565_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg32_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg566_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg372_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg28_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg374_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product310_4_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_4_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Product610_0_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Product610_0_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Product610_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_0_impl_out,
                 X => Delay1No44_out_to_Product610_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Product610_0_impl_parent_implementedSystem_port_1_cast);

SharedReg507_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg507_out;
SharedReg1_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg113_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg113_out;
SharedReg565_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg215_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg215_out;
SharedReg94_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg94_out;
SharedReg113_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg113_out;
SharedReg425_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg425_out;
SharedReg177_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg177_out;
Delay13No30_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_14_cast <= Delay13No30_out;
SharedReg431_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg431_out;
SharedReg557_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg557_out;
   MUX_Product610_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg507_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg113_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg425_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg177_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay13No30_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg431_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg557_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg8_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg113_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg215_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg94_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product610_0_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_0_impl_0_out,
                 Y => Delay1No44_out);

SharedReg571_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg571_out;
SharedReg13_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg31_out;
SharedReg561_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg27_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg27_out;
SharedReg575_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg575_out;
SharedReg33_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg33_out;
SharedReg327_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg327_out;
SharedReg368_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg368_out;
SharedReg576_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg576_out;
SharedReg577_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg577_out;
SharedReg258_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg258_out;
   MUX_Product610_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg571_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg33_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg327_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg368_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg576_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg577_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg258_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg31_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg27_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg575_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product610_0_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_0_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Product610_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_1_impl_out,
                 X => Delay1No46_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast);

SharedReg492_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg492_out;
Delay14No16_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast <= Delay14No16_out;
SharedReg557_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg414_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg414_out;
SharedReg1_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg117_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg117_out;
SharedReg148_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg148_out;
SharedReg565_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg565_out;
SharedReg434_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg434_out;
SharedReg414_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg414_out;
SharedReg500_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg500_out;
SharedReg433_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg433_out;
SharedReg494_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg494_out;
   MUX_Product610_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg492_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay14No16_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg434_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg414_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg500_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg433_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg494_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg414_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg8_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg117_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg148_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product610_1_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_1_impl_0_out,
                 Y => Delay1No46_out);

SharedReg568_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg568_out;
SharedReg577_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg577_out;
SharedReg267_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg267_out;
SharedReg571_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg571_out;
SharedReg13_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg31_out;
SharedReg561_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg565_out;
SharedReg16_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg16_out;
SharedReg566_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg566_out;
SharedReg336_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg336_out;
SharedReg336_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg336_out;
SharedReg311_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg311_out;
   MUX_Product610_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg568_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg577_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg16_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg566_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg336_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg336_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg311_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg267_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg571_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg13_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg31_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product610_1_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_1_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Product610_2_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Product610_2_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Product610_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_2_impl_out,
                 X => Delay1No48_out_to_Product610_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Product610_2_impl_parent_implementedSystem_port_1_cast);

SharedReg4_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg4_out;
SharedReg231_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg231_out;
SharedReg453_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg453_out;
SharedReg451_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg451_out;
SharedReg103_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg103_out;
SharedReg557_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg482_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg482_out;
SharedReg30_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg30_out;
SharedReg2_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg2_out;
SharedReg561_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg123_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg123_out;
SharedReg156_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg156_out;
SharedReg565_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg565_out;
SharedReg420_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg420_out;
SharedReg231_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg231_out;
   MUX_Product610_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg4_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg231_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg123_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg156_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg565_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg420_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg231_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg453_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg451_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg103_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg482_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg30_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg2_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product610_2_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_2_impl_0_out,
                 Y => Delay1No48_out);

SharedReg344_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg344_out;
SharedReg344_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg344_out;
SharedReg293_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg293_out;
SharedReg568_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg568_out;
SharedReg577_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg577_out;
SharedReg275_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg275_out;
SharedReg571_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg571_out;
SharedReg20_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg565_out;
SharedReg27_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg27_out;
SharedReg566_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg566_out;
   MUX_Product610_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg344_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg344_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg564_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg565_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg27_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg566_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg293_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg568_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg577_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg275_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg571_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg20_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg26_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product610_2_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_2_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Product610_3_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Product610_3_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Product610_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_3_impl_out,
                 X => Delay1No50_out_to_Product610_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Product610_3_impl_parent_implementedSystem_port_1_cast);

SharedReg478_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg478_out;
SharedReg237_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg237_out;
SharedReg400_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg400_out;
SharedReg236_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg236_out;
SharedReg60_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg60_out;
SharedReg132_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg132_out;
SharedReg460_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg460_out;
SharedReg111_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg111_out;
SharedReg557_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg476_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg476_out;
SharedReg30_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg30_out;
SharedReg2_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg2_out;
SharedReg561_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg130_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg130_out;
SharedReg163_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg163_out;
   MUX_Product610_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg478_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg237_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg30_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg2_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg130_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg163_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg400_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg236_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg60_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg132_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg460_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg111_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg476_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product610_3_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_3_impl_0_out,
                 Y => Delay1No50_out);

SharedReg574_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg574_out;
SharedReg16_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg566_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg566_out;
SharedReg567_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg567_out;
SharedReg284_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg284_out;
SharedReg300_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg300_out;
SharedReg568_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg568_out;
SharedReg577_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg577_out;
SharedReg289_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg289_out;
SharedReg571_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg571_out;
SharedReg20_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg564_out;
   MUX_Product610_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg574_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg26_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg564_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg566_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg567_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg284_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg300_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg568_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg577_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg289_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg571_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product610_3_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_3_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Product610_4_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Product610_4_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Product610_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_4_impl_out,
                 X => Delay1No52_out_to_Product610_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Product610_4_impl_parent_implementedSystem_port_1_cast);

SharedReg561_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg563_out;
SharedReg243_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg243_out;
SharedReg477_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg477_out;
SharedReg209_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg209_out;
SharedReg443_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg443_out;
SharedReg465_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg465_out;
SharedReg439_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg439_out;
SharedReg373_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg373_out;
SharedReg362_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg362_out;
SharedReg213_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg213_out;
SharedReg557_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg557_out;
SharedReg209_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg209_out;
SharedReg1_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1_out;
SharedReg2_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg2_out;
   MUX_Product610_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg362_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg213_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg557_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg209_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg2_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg563_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg243_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg477_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg209_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg443_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg465_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg439_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg373_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product610_4_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_4_impl_0_out,
                 Y => Delay1No52_out);

SharedReg561_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg9_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg9_out;
SharedReg21_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg21_out;
SharedReg575_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg575_out;
SharedReg359_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg359_out;
SharedReg5_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg5_out;
SharedReg374_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg374_out;
SharedReg375_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg375_out;
SharedReg577_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg577_out;
Delay131No4_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_13_cast <= Delay131No4_out;
SharedReg571_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg571_out;
SharedReg13_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg13_out;
SharedReg26_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg26_out;
   MUX_Product610_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg375_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg577_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay131No4_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg571_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg13_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg26_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg563_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg9_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg21_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg575_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg359_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg5_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg374_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product610_4_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_4_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Product810_0_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Product810_0_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Product810_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_0_impl_out,
                 X => Delay1No54_out_to_Product810_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Product810_0_impl_parent_implementedSystem_port_1_cast);

SharedReg519_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg519_out;
SharedReg30_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg30_out;
SharedReg2_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg561_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg113_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg113_out;
SharedReg141_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg141_out;
SharedReg565_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg408_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg408_out;
SharedReg507_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg507_out;
SharedReg528_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg528_out;
SharedReg407_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg407_out;
SharedReg522_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg522_out;
SharedReg329_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg329_out;
SharedReg527_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg527_out;
SharedReg557_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg557_out;
   MUX_Product810_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg519_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg528_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg407_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg522_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg329_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg527_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg557_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg2_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg113_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg141_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg408_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg507_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product810_0_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_0_impl_0_out,
                 Y => Delay1No54_out);

SharedReg571_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg571_out;
SharedReg20_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg16_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg16_out;
SharedReg566_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg566_out;
SharedReg367_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg367_out;
SharedReg367_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg367_out;
SharedReg328_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg328_out;
SharedReg24_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg24_out;
SharedReg569_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg569_out;
SharedReg334_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg334_out;
   MUX_Product810_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg571_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg367_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg367_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg328_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg24_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg569_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg334_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg26_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg16_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg566_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product810_0_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_0_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Product810_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_1_impl_out,
                 X => Delay1No56_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast);

SharedReg501_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg501_out;
SharedReg499_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg499_out;
SharedReg557_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg490_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg490_out;
SharedReg30_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg30_out;
SharedReg2_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg2_out;
SharedReg561_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg148_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg148_out;
SharedReg183_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg183_out;
SharedReg565_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg565_out;
SharedReg415_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg415_out;
SharedReg433_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg433_out;
SharedReg414_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg414_out;
SharedReg336_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg336_out;
SharedReg149_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg149_out;
   MUX_Product810_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg501_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg499_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg415_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg433_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg414_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg336_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg149_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg490_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg30_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg2_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg148_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg183_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product810_1_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_1_impl_0_out,
                 Y => Delay1No56_out);

SharedReg568_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg568_out;
SharedReg569_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg569_out;
SharedReg342_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg342_out;
SharedReg571_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg571_out;
SharedReg20_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg565_out;
SharedReg27_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg27_out;
SharedReg566_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg566_out;
SharedReg567_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg567_out;
SharedReg28_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg28_out;
SharedReg29_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg29_out;
   MUX_Product810_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg568_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg569_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg27_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg566_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg567_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg28_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg29_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg342_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg571_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg26_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product810_1_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_1_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Product810_2_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Product810_2_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Product810_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_2_impl_out,
                 X => Delay1No58_out_to_Product810_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Product810_2_impl_parent_implementedSystem_port_1_cast);

SharedReg565_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg344_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg344_out;
SharedReg124_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg124_out;
SharedReg484_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg484_out;
SharedReg191_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg191_out;
SharedReg557_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg392_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg392_out;
SharedReg1_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg191_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg191_out;
SharedReg191_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg191_out;
SharedReg565_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg565_out;
SharedReg124_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg124_out;
SharedReg449_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg449_out;
   MUX_Product810_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg344_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg191_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg191_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg565_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg124_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg449_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg124_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg484_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg191_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg392_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg8_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product810_2_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_2_impl_0_out,
                 Y => Delay1No58_out);

SharedReg565_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg28_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg28_out;
SharedReg29_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg29_out;
SharedReg568_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg568_out;
SharedReg569_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg569_out;
SharedReg274_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg274_out;
SharedReg571_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg571_out;
SharedReg20_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg565_out;
SharedReg16_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg16_out;
SharedReg566_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg566_out;
   MUX_Product810_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg28_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg564_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg565_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg16_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg566_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg29_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg568_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg569_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg274_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg571_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg20_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg26_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product810_2_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_2_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Product810_3_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Product810_3_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Product810_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_3_impl_out,
                 X => Delay1No60_out_to_Product810_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Product810_3_impl_parent_implementedSystem_port_1_cast);

SharedReg561_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg401_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg401_out;
SharedReg236_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg236_out;
SharedReg4_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg4_out;
SharedReg105_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg105_out;
SharedReg462_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg462_out;
SharedReg472_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg472_out;
SharedReg236_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg236_out;
SharedReg557_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg70_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg70_out;
SharedReg1_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg199_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg199_out;
SharedReg199_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg199_out;
   MUX_Product810_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg401_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg8_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg199_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg199_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg236_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg4_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg105_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg462_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg472_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg236_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg70_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product810_3_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_3_impl_0_out,
                 Y => Delay1No60_out);

SharedReg561_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg27_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg27_out;
SharedReg566_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg566_out;
SharedReg299_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg299_out;
SharedReg299_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg299_out;
SharedReg285_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg285_out;
SharedReg568_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg568_out;
SharedReg569_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg569_out;
Delay125No3_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_9_cast <= Delay125No3_out;
SharedReg571_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg571_out;
SharedReg20_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg564_out;
   MUX_Product810_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg26_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg564_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg566_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg299_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg299_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg285_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg568_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg569_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay125No3_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg571_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product810_3_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_3_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Product810_4_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Product810_4_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Product810_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_4_impl_out,
                 X => Delay1No62_out_to_Product810_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Product810_4_impl_parent_implementedSystem_port_1_cast);

SharedReg561_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg137_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg137_out;
SharedReg513_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg513_out;
SharedReg565_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg565_out;
SharedReg243_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg243_out;
SharedReg535_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg535_out;
SharedReg469_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg469_out;
SharedReg464_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg464_out;
SharedReg361_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg361_out;
SharedReg173_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg173_out;
SharedReg467_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg467_out;
SharedReg557_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg557_out;
SharedReg243_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg243_out;
SharedReg30_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg30_out;
SharedReg8_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg8_out;
   MUX_Product810_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg173_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg467_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg557_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg243_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg30_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg8_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg137_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg513_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg565_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg243_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg535_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg469_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg464_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg361_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product810_4_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_4_impl_0_out,
                 Y => Delay1No62_out);

SharedReg561_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg565_out;
SharedReg27_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg27_out;
SharedReg566_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg566_out;
SharedReg33_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg33_out;
SharedReg360_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg360_out;
SharedReg373_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg373_out;
SharedReg576_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg576_out;
SharedReg577_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg577_out;
SharedReg366_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg366_out;
SharedReg571_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg571_out;
SharedReg20_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg26_out;
   MUX_Product810_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg576_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg577_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg366_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg571_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg20_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg26_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg563_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg565_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg27_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg566_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg33_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg360_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg373_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product810_4_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_4_impl_1_out,
                 Y => Delay1No63_out);
   Inv_11_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_0_IEEE,
                 X => Delay1No64_out);
Inv_11_0 <= Inv_11_0_IEEE;

SharedReg40_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_1_cast <= SharedReg40_out;
SharedReg48_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_2_cast <= SharedReg48_out;
SharedReg54_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_3_cast <= SharedReg54_out;
SharedReg60_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_4_cast <= SharedReg60_out;
SharedReg64_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_5_cast <= SharedReg64_out;
   MUX_Inv_11_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg40_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg48_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg54_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg64_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_11_0_0_LUT_out,
                 oMux => MUX_Inv_11_0_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_11_0_0_out,
                 Y => Delay1No64_out);
   Inv_12_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_0_IEEE,
                 X => Delay1No65_out);
Inv_12_0 <= Inv_12_0_IEEE;

SharedReg40_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_1_cast <= SharedReg40_out;
SharedReg48_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_2_cast <= SharedReg48_out;
SharedReg54_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_3_cast <= SharedReg54_out;
SharedReg60_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_4_cast <= SharedReg60_out;
SharedReg70_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_5_cast <= SharedReg70_out;
   MUX_Inv_12_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg40_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg48_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg54_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg70_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_12_0_0_LUT_out,
                 oMux => MUX_Inv_12_0_0_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_12_0_0_out,
                 Y => Delay1No65_out);
   Inv_13_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_0_IEEE,
                 X => Delay1No66_out);
Inv_13_0 <= Inv_13_0_IEEE;

SharedReg113_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_1_cast <= SharedReg113_out;
SharedReg117_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
SharedReg123_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_3_cast <= SharedReg123_out;
SharedReg130_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_4_cast <= SharedReg130_out;
SharedReg137_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_5_cast <= SharedReg137_out;
   MUX_Inv_13_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg113_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg123_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg130_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg137_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_13_0_0_LUT_out,
                 oMux => MUX_Inv_13_0_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_13_0_0_out,
                 Y => Delay1No66_out);
   Inv_21_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_0_IEEE,
                 X => Delay1No67_out);
Inv_21_0 <= Inv_21_0_IEEE;

SharedReg141_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_1_cast <= SharedReg141_out;
SharedReg148_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_2_cast <= SharedReg148_out;
SharedReg156_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_3_cast <= SharedReg156_out;
SharedReg163_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_4_cast <= SharedReg163_out;
SharedReg169_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_5_cast <= SharedReg169_out;
   MUX_Inv_21_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg141_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg148_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg156_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg163_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg169_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_21_0_0_LUT_out,
                 oMux => MUX_Inv_21_0_0_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_21_0_0_out,
                 Y => Delay1No67_out);
   Inv_22_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_0_IEEE,
                 X => Delay1No68_out);
Inv_22_0 <= Inv_22_0_IEEE;

SharedReg89_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_1_cast <= SharedReg89_out;
SharedReg95_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_2_cast <= SharedReg95_out;
SharedReg54_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_3_cast <= SharedReg54_out;
SharedReg60_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_4_cast <= SharedReg60_out;
SharedReg64_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_5_cast <= SharedReg64_out;
   MUX_Inv_22_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg89_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg95_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg54_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg64_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_22_0_0_LUT_out,
                 oMux => MUX_Inv_22_0_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_22_0_0_out,
                 Y => Delay1No68_out);
   Inv_23_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_0_IEEE,
                 X => Delay1No69_out);
Inv_23_0 <= Inv_23_0_IEEE;

SharedReg113_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_1_cast <= SharedReg113_out;
SharedReg117_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
SharedReg99_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_3_cast <= SharedReg99_out;
SharedReg105_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_4_cast <= SharedReg105_out;
SharedReg137_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_5_cast <= SharedReg137_out;
   MUX_Inv_23_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg113_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg99_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg137_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_23_0_0_LUT_out,
                 oMux => MUX_Inv_23_0_0_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_23_0_0_out,
                 Y => Delay1No69_out);
   Inv_31_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_0_IEEE,
                 X => Delay1No70_out);
Inv_31_0 <= Inv_31_0_IEEE;

SharedReg175_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_1_cast <= SharedReg175_out;
SharedReg183_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_2_cast <= SharedReg183_out;
SharedReg191_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_3_cast <= SharedReg191_out;
SharedReg199_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_4_cast <= SharedReg199_out;
SharedReg209_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_5_cast <= SharedReg209_out;
   MUX_Inv_31_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg175_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg183_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg191_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg199_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg209_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_31_0_0_LUT_out,
                 oMux => MUX_Inv_31_0_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_31_0_0_out,
                 Y => Delay1No70_out);
   Inv_32_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_0_IEEE,
                 X => Delay1No71_out);
Inv_32_0 <= Inv_32_0_IEEE;

SharedReg89_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_1_cast <= SharedReg89_out;
SharedReg95_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_2_cast <= SharedReg95_out;
SharedReg99_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_3_cast <= SharedReg99_out;
SharedReg105_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_4_cast <= SharedReg105_out;
SharedReg137_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_5_cast <= SharedReg137_out;
   MUX_Inv_32_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg89_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg95_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg99_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg137_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_32_0_0_LUT_out,
                 oMux => MUX_Inv_32_0_0_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_32_0_0_out,
                 Y => Delay1No71_out);
   Inv_33_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_0_IEEE,
                 X => Delay1No72_out);
Inv_33_0 <= Inv_33_0_IEEE;

SharedReg215_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_1_cast <= SharedReg215_out;
SharedReg223_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_2_cast <= SharedReg223_out;
SharedReg231_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_3_cast <= SharedReg231_out;
SharedReg236_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_4_cast <= SharedReg236_out;
SharedReg243_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_5_cast <= SharedReg243_out;
   MUX_Inv_33_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg215_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg223_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg231_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg236_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg243_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_33_0_0_LUT_out,
                 oMux => MUX_Inv_33_0_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_33_0_0_out,
                 Y => Delay1No72_out);
   Inv_41_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_0_IEEE,
                 X => Delay1No73_out);
Inv_41_0 <= Inv_41_0_IEEE;

SharedReg130_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_1_cast <= SharedReg130_out;
SharedReg113_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_2_cast <= SharedReg113_out;
SharedReg117_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_3_cast <= SharedReg117_out;
SharedReg123_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_4_cast <= SharedReg123_out;
SharedReg169_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_5_cast <= SharedReg169_out;
   MUX_Inv_41_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg130_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg113_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg117_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg123_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg169_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_41_0_0_LUT_out,
                 oMux => MUX_Inv_41_0_0_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_41_0_0_out,
                 Y => Delay1No73_out);
   Inv_42_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_0_IEEE,
                 X => Delay1No74_out);
Inv_42_0 <= Inv_42_0_IEEE;

SharedReg40_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_1_cast <= SharedReg40_out;
SharedReg48_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_2_cast <= SharedReg48_out;
SharedReg76_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_3_cast <= SharedReg76_out;
SharedReg82_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_4_cast <= SharedReg82_out;
SharedReg70_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_5_cast <= SharedReg70_out;
   MUX_Inv_42_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg40_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg48_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg76_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg82_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg70_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_42_0_0_LUT_out,
                 oMux => MUX_Inv_42_0_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_42_0_0_out,
                 Y => Delay1No74_out);
   Inv_43_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_0_IEEE,
                 X => Delay1No75_out);
Inv_43_0 <= Inv_43_0_IEEE;

SharedReg89_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_1_cast <= SharedReg89_out;
SharedReg95_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_2_cast <= SharedReg95_out;
SharedReg99_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_3_cast <= SharedReg99_out;
SharedReg105_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_4_cast <= SharedReg105_out;
SharedReg64_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_5_cast <= SharedReg64_out;
   MUX_Inv_43_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg89_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg95_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg99_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg64_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_43_0_0_LUT_out,
                 oMux => MUX_Inv_43_0_0_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_43_0_0_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Add30_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_0_impl_out,
                 X => Delay1No76_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast);

SharedReg141_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg141_out;
Delay25No_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast <= Delay25No_out;
SharedReg141_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg141_out;
SharedReg512_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg512_out;
SharedReg175_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg175_out;
SharedReg182_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg182_out;
SharedReg45_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg45_out;
SharedReg144_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg144_out;
SharedReg178_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg178_out;
SharedReg146_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg146_out;
SharedReg47_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg47_out;
SharedReg531_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg531_out;
SharedReg407_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg407_out;
SharedReg141_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg141_out;
SharedReg221_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg221_out;
SharedReg175_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg175_out;
   MUX_Add30_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg141_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay25No_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg47_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg531_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg407_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg141_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg221_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg175_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg141_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg512_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg182_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg45_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg144_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg178_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg146_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add30_0_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_0_impl_0_out,
                 Y => Delay1No76_out);

SharedReg217_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg217_out;
SharedReg546_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg546_out;
SharedReg332_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg332_out;
SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg545_out;
SharedReg430_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg430_out;
SharedReg367_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg367_out;
SharedReg251_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg251_out;
SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg545_out;
SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg545_out;
SharedReg251_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg251_out;
SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg545_out;
SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg545_out;
SharedReg507_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg507_out;
SharedReg216_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg216_out;
SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg545_out;
SharedReg215_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg215_out;
   MUX_Add30_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg217_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg546_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg507_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg216_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg215_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg332_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg430_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg367_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg251_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg545_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg251_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add30_0_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_0_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Add30_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_1_impl_out,
                 X => Delay1No78_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast);

SharedReg113_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg113_out;
Delay59No_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast <= Delay59No_out;
SharedReg534_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg534_out;
SharedReg117_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg117_out;
SharedReg497_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg497_out;
SharedReg148_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg148_out;
SharedReg496_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg496_out;
SharedReg183_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg183_out;
SharedReg155_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg155_out;
SharedReg410_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg410_out;
SharedReg120_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg120_out;
SharedReg151_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg151_out;
SharedReg121_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg121_out;
SharedReg382_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg382_out;
SharedReg505_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg505_out;
SharedReg433_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg433_out;
   MUX_Add30_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg113_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay59No_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg120_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg151_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg121_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg382_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg505_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg433_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg534_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg117_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg497_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg148_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg496_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg183_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg155_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg410_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add30_1_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_1_impl_0_out,
                 Y => Delay1No78_out);

SharedReg114_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg114_out;
SharedReg545_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg545_out;
SharedReg328_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg328_out;
SharedReg185_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg185_out;
SharedReg336_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg336_out;
SharedReg315_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg315_out;
SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg547_out;
SharedReg228_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg228_out;
SharedReg336_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg336_out;
SharedReg326_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg326_out;
SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg547_out;
SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg547_out;
SharedReg259_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg259_out;
SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg547_out;
SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg547_out;
SharedReg414_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg414_out;
   MUX_Add30_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg114_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg545_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg259_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg414_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg328_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg185_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg336_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg315_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg547_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg228_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg336_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg326_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add30_1_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_1_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Add30_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_2_impl_out,
                 X => Delay1No80_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast);

SharedReg414_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg414_out;
SharedReg498_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg498_out;
SharedReg48_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg48_out;
SharedReg95_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg95_out;
SharedReg126_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg126_out;
Delay81No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_6_cast <= Delay81No1_out;
SharedReg123_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg123_out;
SharedReg162_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg162_out;
SharedReg156_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg156_out;
SharedReg487_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg487_out;
SharedReg156_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg156_out;
SharedReg128_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg128_out;
SharedReg416_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg416_out;
SharedReg503_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg503_out;
SharedReg159_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg159_out;
SharedReg104_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg104_out;
   MUX_Add30_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg414_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg498_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg156_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg128_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg416_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg503_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg159_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg104_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg48_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg95_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg126_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay81No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg123_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg162_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg156_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg487_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add30_2_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_2_impl_0_out,
                 Y => Delay1No80_out);

SharedReg496_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg496_out;
SharedReg338_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg338_out;
SharedReg49_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg49_out;
SharedReg96_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg96_out;
SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg549_out;
SharedReg311_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg311_out;
SharedReg78_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg78_out;
SharedReg276_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg276_out;
SharedReg349_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg349_out;
SharedReg550_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg550_out;
SharedReg195_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg195_out;
SharedReg344_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg344_out;
SharedReg309_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg309_out;
SharedReg550_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg550_out;
SharedReg550_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg550_out;
SharedReg268_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg268_out;
   MUX_Add30_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg496_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg338_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg195_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg344_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg309_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg550_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg550_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg268_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg49_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg96_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg311_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg78_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg276_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg349_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg550_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add30_2_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_2_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Add30_3_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Add30_3_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Add30_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_3_impl_out,
                 X => Delay1No82_out_to_Add30_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Add30_3_impl_parent_implementedSystem_port_1_cast);

SharedReg489_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg489_out;
Delay90No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_2_cast <= Delay90No2_out;
Delay32No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_3_cast <= Delay32No2_out;
SharedReg419_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg419_out;
Delay111No3_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_5_cast <= Delay111No3_out;
SharedReg54_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg54_out;
SharedReg99_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg99_out;
SharedReg166_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg166_out;
Delay81No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_9_cast <= Delay81No2_out;
SharedReg163_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg163_out;
SharedReg207_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg207_out;
SharedReg163_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg163_out;
SharedReg475_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg475_out;
SharedReg163_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg163_out;
SharedReg168_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg168_out;
SharedReg422_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg422_out;
   MUX_Add30_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg489_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay90No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg207_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg163_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg475_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg163_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg168_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg422_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => Delay32No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg419_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay111No3_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg54_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg99_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg166_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay81No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg163_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add30_3_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_3_impl_0_out,
                 Y => Delay1No82_out);

SharedReg340_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg340_out;
SharedReg280_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg280_out;
SharedReg291_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg291_out;
SharedReg455_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg455_out;
SharedReg303_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg303_out;
SharedReg415_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg415_out;
SharedReg491_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg491_out;
SharedReg549_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg549_out;
SharedReg346_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg346_out;
SharedReg61_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg61_out;
SharedReg353_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg353_out;
SharedReg305_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg305_out;
SharedReg551_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg551_out;
SharedReg204_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg204_out;
SharedReg299_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg299_out;
SharedReg291_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg291_out;
   MUX_Add30_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg340_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg280_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg353_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg305_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg551_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg204_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg299_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg291_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg291_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg455_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg303_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg415_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg491_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg549_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg346_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg61_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add30_3_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_3_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Add30_4_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Add30_4_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Add30_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_4_impl_out,
                 X => Delay1No84_out_to_Add30_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Add30_4_impl_parent_implementedSystem_port_1_cast);

SharedReg396_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg396_out;
SharedReg202_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg202_out;
SharedReg112_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg112_out;
SharedReg87_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg87_out;
Delay90No3_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_5_cast <= Delay90No3_out;
SharedReg400_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg400_out;
SharedReg130_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg130_out;
SharedReg463_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg463_out;
SharedReg199_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg199_out;
SharedReg473_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg473_out;
SharedReg481_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg481_out;
SharedReg242_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg242_out;
SharedReg458_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg458_out;
SharedReg476_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg476_out;
SharedReg_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg_out;
SharedReg63_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg63_out;
   MUX_Add30_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg396_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg202_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg481_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg242_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg458_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg476_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg63_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg112_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg87_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay90No3_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg400_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg130_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg463_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg199_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg473_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add30_4_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_4_impl_0_out,
                 Y => Delay1No84_out);

SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg551_out;
SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg551_out;
SharedReg276_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg276_out;
SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg551_out;
SharedReg356_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg356_out;
SharedReg458_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg458_out;
SharedReg200_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg200_out;
SharedReg354_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg354_out;
SharedReg236_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg236_out;
SharedReg400_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg400_out;
SharedReg550_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg550_out;
SharedReg353_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg353_out;
SharedReg304_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg304_out;
SharedReg441_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg441_out;
SharedReg476_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg476_out;
SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg551_out;
   MUX_Add30_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg550_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg353_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg304_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg441_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg476_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg276_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg356_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg458_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg200_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg354_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg236_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg400_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add30_4_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_4_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Add110_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_2_impl_out,
                 X => Delay1No86_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast);

SharedReg389_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg389_out;
SharedReg486_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg486_out;
SharedReg231_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg231_out;
SharedReg99_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg99_out;
SharedReg456_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg456_out;
SharedReg156_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg156_out;
SharedReg452_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg452_out;
Delay59No2_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_8_cast <= Delay59No2_out;
SharedReg235_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg235_out;
SharedReg449_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg449_out;
SharedReg399_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg399_out;
SharedReg_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg_out;
SharedReg81_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg81_out;
SharedReg198_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg198_out;
SharedReg127_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg127_out;
SharedReg76_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg76_out;
   MUX_Add110_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg389_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg486_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg399_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg81_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg198_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg127_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg76_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg231_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg99_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg456_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg156_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg452_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay59No2_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg235_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg449_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add110_2_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_2_impl_0_out,
                 Y => Delay1No86_out);

SharedReg550_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg550_out;
SharedReg550_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg550_out;
SharedReg419_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg419_out;
SharedReg157_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg157_out;
SharedReg346_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg346_out;
SharedReg191_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg191_out;
SharedReg231_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg231_out;
SharedReg547_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg547_out;
SharedReg276_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg276_out;
SharedReg296_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg296_out;
SharedReg552_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg552_out;
SharedReg392_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg392_out;
SharedReg550_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg550_out;
SharedReg291_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg291_out;
SharedReg268_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg268_out;
SharedReg54_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg54_out;
   MUX_Add110_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg550_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg550_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg552_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg392_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg550_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg291_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg268_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg54_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg419_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg157_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg346_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg191_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg231_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg547_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg276_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg296_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add110_2_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_2_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Add110_4_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Add110_4_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Add110_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_4_impl_out,
                 X => Delay1No88_out_to_Add110_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Add110_4_impl_parent_implementedSystem_port_1_cast);

SharedReg206_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg206_out;
SharedReg135_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg135_out;
SharedReg82_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg82_out;
SharedReg163_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg163_out;
SharedReg212_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg212_out;
SharedReg130_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg130_out;
SharedReg488_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg488_out;
SharedReg405_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg405_out;
SharedReg61_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg61_out;
SharedReg88_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg88_out;
SharedReg476_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg476_out;
Delay88No3_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_12_cast <= Delay88No3_out;
Delay35No3_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_13_cast <= Delay35No3_out;
SharedReg537_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg537_out;
SharedReg36_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg36_out;
SharedReg19_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg19_out;
   MUX_Add110_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg206_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg135_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg476_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay88No3_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay35No3_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg537_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg36_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg19_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg82_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg163_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg212_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg130_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg488_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg405_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg61_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg88_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add110_4_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_4_impl_0_out,
                 Y => Delay1No88_out);

SharedReg283_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg283_out;
SharedReg276_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg276_out;
SharedReg60_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg60_out;
SharedReg199_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg199_out;
SharedReg551_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg551_out;
SharedReg163_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg163_out;
SharedReg551_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg551_out;
SharedReg551_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg551_out;
SharedReg60_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg60_out;
SharedReg548_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg548_out;
SharedReg440_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg440_out;
SharedReg355_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg355_out;
SharedReg283_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg283_out;
SharedReg137_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg137_out;
SharedReg70_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg70_out;
SharedReg70_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg70_out;
   MUX_Add110_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg283_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg276_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg440_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg355_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg283_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg137_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg70_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg70_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg60_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg199_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg551_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg163_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg551_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg551_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg60_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg548_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add110_4_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_4_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Add101_1_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Add101_1_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Add101_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add101_1_impl_out,
                 X => Delay1No90_out_to_Add101_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Add101_1_impl_parent_implementedSystem_port_1_cast);

SharedReg117_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg188_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg188_out;
SharedReg148_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg148_out;
SharedReg493_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg493_out;
SharedReg391_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg391_out;
SharedReg229_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg229_out;
SharedReg414_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg414_out;
SharedReg390_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg390_out;
SharedReg_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg_out;
SharedReg53_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg53_out;
SharedReg190_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg190_out;
SharedReg154_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg154_out;
SharedReg48_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg48_out;
SharedReg183_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg183_out;
Delay111No1_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_15_cast <= Delay111No1_out;
SharedReg117_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg117_out;
   MUX_Add101_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg188_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg190_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg154_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg48_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg183_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay111No1_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg117_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg148_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg493_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg391_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg229_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg414_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg390_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg53_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add101_1_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_1_impl_0_out,
                 Y => Delay1No90_out);

SharedReg184_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg184_out;
SharedReg547_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg547_out;
SharedReg183_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg183_out;
SharedReg223_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg223_out;
SharedReg545_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg545_out;
SharedReg268_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg268_out;
SharedReg314_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg314_out;
Delay2No132_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_8_cast <= Delay2No132_out;
SharedReg385_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg385_out;
SharedReg547_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg547_out;
SharedReg309_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg309_out;
SharedReg259_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg259_out;
SharedReg95_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg95_out;
SharedReg223_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg223_out;
SharedReg340_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg340_out;
SharedReg148_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg148_out;
   MUX_Add101_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg184_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg547_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg309_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg259_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg95_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg223_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg340_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg148_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg183_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg223_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg545_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg268_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg314_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay2No132_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg385_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg547_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add101_1_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_1_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Add121_4_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Add121_4_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Add121_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_4_impl_out,
                 X => Delay1No92_out_to_Add121_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Add121_4_impl_parent_implementedSystem_port_1_cast);

SharedReg514_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg514_out;
SharedReg209_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg209_out;
SharedReg74_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg74_out;
SharedReg67_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg67_out;
Delay43No4_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_5_cast <= Delay43No4_out;
SharedReg73_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg73_out;
SharedReg480_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg480_out;
SharedReg544_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg544_out;
SharedReg542_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg542_out;
SharedReg513_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg513_out;
SharedReg209_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg209_out;
SharedReg69_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg69_out;
SharedReg459_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg459_out;
SharedReg469_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg469_out;
Delay84No4_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_15_cast <= Delay84No4_out;
SharedReg543_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg543_out;
   MUX_Add121_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg514_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg209_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg209_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg69_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg459_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg469_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay84No4_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg543_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg74_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg67_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay43No4_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg73_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg480_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg544_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg542_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg513_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add121_4_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_4_impl_0_out,
                 Y => Delay1No92_out);

SharedReg553_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg553_out;
SharedReg445_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg445_out;
SharedReg353_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg353_out;
SharedReg353_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg353_out;
SharedReg360_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg360_out;
SharedReg550_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg550_out;
SharedReg318_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg318_out;
SharedReg321_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg321_out;
SharedReg550_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg550_out;
SharedReg516_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg516_out;
SharedReg250_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg250_out;
SharedReg550_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg550_out;
SharedReg64_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg64_out;
SharedReg171_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg171_out;
SharedReg376_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg376_out;
SharedReg318_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg318_out;
   MUX_Add121_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg553_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg445_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg250_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg550_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg64_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg171_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg376_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg318_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg353_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg360_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg550_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg318_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg321_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg550_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg516_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add121_4_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_4_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Add141_0_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Add141_0_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Add141_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add141_0_impl_out,
                 X => Delay1No94_out_to_Add141_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Add141_0_impl_parent_implementedSystem_port_1_cast);

SharedReg521_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg521_out;
Delay84No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_2_cast <= Delay84No_out;
SharedReg532_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg532_out;
SharedReg407_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg407_out;
SharedReg384_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg384_out;
SharedReg_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg_out;
Delay11No40_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_7_cast <= Delay11No40_out;
SharedReg525_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg525_out;
Delay21No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_9_cast <= Delay21No_out;
SharedReg89_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg89_out;
SharedReg215_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg215_out;
Delay111No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_12_cast <= Delay111No_out;
SharedReg141_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg141_out;
SharedReg147_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg147_out;
SharedReg146_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg146_out;
SharedReg91_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg91_out;
   MUX_Add141_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg521_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay84No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg215_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay111No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg141_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg147_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg146_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg91_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg532_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg407_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg384_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay11No40_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg525_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay21No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg89_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add141_0_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_0_impl_0_out,
                 Y => Delay1No94_out);

SharedReg425_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg425_out;
SharedReg371_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg371_out;
SharedReg367_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg367_out;
SharedReg331_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg331_out;
SharedReg548_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg548_out;
SharedReg527_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg527_out;
SharedReg545_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg545_out;
SharedReg326_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg326_out;
SharedReg251_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg251_out;
SharedReg113_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg113_out;
SharedReg425_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg425_out;
SharedReg371_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg371_out;
SharedReg175_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg175_out;
SharedReg545_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg545_out;
Delay3No65_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_15_cast <= Delay3No65_out;
SharedReg40_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg40_out;
   MUX_Add141_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg425_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg371_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg425_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg371_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg175_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg545_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay3No65_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg40_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg367_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg331_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg548_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg527_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg545_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg326_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg251_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg113_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add141_0_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_0_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Add151_2_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Add151_2_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Add151_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add151_2_impl_out,
                 X => Delay1No96_out_to_Add151_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Add151_2_impl_parent_implementedSystem_port_1_cast);

SharedReg122_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg122_out;
SharedReg121_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg121_out;
SharedReg50_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg50_out;
SharedReg383_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg383_out;
SharedReg197_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg197_out;
Delay88No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_6_cast <= Delay88No1_out;
Delay35No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_7_cast <= Delay35No1_out;
Delay84No2_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_8_cast <= Delay84No2_out;
SharedReg36_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg36_out;
SharedReg19_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg19_out;
Delay43No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_11_cast <= Delay43No1_out;
SharedReg418_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg418_out;
SharedReg382_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg382_out;
SharedReg506_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg506_out;
Delay90No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_15_cast <= Delay90No1_out;
Delay32No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_16_cast <= Delay32No1_out;
   MUX_Add151_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg122_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg121_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay43No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg418_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg382_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg506_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay90No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay32No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg50_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg383_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg197_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay88No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay35No1_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay84No2_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg36_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg19_out_to_MUX_Add151_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add151_2_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add151_2_impl_0_out,
                 Y => Delay1No96_out);

SharedReg547_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg547_out;
SharedReg549_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg549_out;
SharedReg377_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg377_out;
SharedReg546_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg546_out;
SharedReg547_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg547_out;
SharedReg339_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg339_out;
SharedReg268_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg268_out;
SharedReg348_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg348_out;
SharedReg76_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg76_out;
SharedReg76_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg76_out;
SharedReg260_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg260_out;
SharedReg311_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg311_out;
SharedReg547_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg547_out;
SharedReg371_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg371_out;
SharedReg271_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg271_out;
SharedReg309_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg309_out;
   MUX_Add151_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg547_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg549_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg260_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg311_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg547_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg371_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg271_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg309_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg377_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg546_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg547_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg339_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg268_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg348_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg76_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg76_out_to_MUX_Add151_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add151_2_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add151_2_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Add151_3_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Add151_3_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Add151_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add151_3_impl_out,
                 X => Delay1No98_out_to_Add151_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Add151_3_impl_parent_implementedSystem_port_1_cast);

SharedReg156_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg156_out;
Delay111No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_2_cast <= Delay111No2_out;
SharedReg99_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg99_out;
Delay19No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_4_cast <= Delay19No2_out;
SharedReg480_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg480_out;
SharedReg78_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg78_out;
Delay16No17_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_7_cast <= Delay16No17_out;
SharedReg241_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg241_out;
SharedReg457_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg457_out;
Delay35No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_10_cast <= Delay35No2_out;
Delay84No3_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_11_cast <= Delay84No3_out;
SharedReg36_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg36_out;
SharedReg19_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg19_out;
Delay43No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_14_cast <= Delay43No2_out;
Delay67No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_15_cast <= Delay67No2_out;
SharedReg389_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg389_out;
   MUX_Add151_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg156_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay111No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay84No3_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg36_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg19_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay43No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay67No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg389_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg99_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay19No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg480_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg78_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay16No17_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg241_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg457_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay35No2_out_to_MUX_Add151_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add151_3_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add151_3_impl_0_out,
                 Y => Delay1No98_out);

SharedReg191_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg191_out;
SharedReg348_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg348_out;
SharedReg123_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg123_out;
SharedReg550_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg550_out;
SharedReg550_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg550_out;
SharedReg76_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg76_out;
SharedReg546_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg546_out;
SharedReg550_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg550_out;
SharedReg279_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg279_out;
SharedReg291_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg291_out;
SharedReg356_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg356_out;
SharedReg82_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg82_out;
SharedReg82_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg82_out;
SharedReg269_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg269_out;
SharedReg293_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg293_out;
SharedReg550_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg550_out;
   MUX_Add151_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg191_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg348_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg356_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg82_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg82_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg269_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg293_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg550_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg123_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg550_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg550_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg76_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg546_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg550_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg279_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg291_out_to_MUX_Add151_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add151_3_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add151_3_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Add16_4_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Add16_4_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Add16_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add16_4_impl_out,
                 X => Delay1No100_out_to_Add16_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Add16_4_impl_parent_implementedSystem_port_1_cast);

SharedReg208_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg208_out;
Delay67No3_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_2_cast <= Delay67No3_out;
SharedReg87_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg87_out;
Delay80No3_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_4_cast <= Delay80No3_out;
SharedReg539_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg539_out;
SharedReg406_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg406_out;
SharedReg458_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg458_out;
SharedReg64_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg64_out;
SharedReg105_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg105_out;
SharedReg130_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg130_out;
Delay19No4_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_11_cast <= Delay19No4_out;
Delay81No3_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_12_cast <= Delay81No3_out;
SharedReg243_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg243_out;
SharedReg249_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg249_out;
SharedReg74_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg74_out;
SharedReg209_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg209_out;
   MUX_Add16_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg208_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay67No3_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay19No4_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay81No3_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg243_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg249_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg74_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg209_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg87_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay80No3_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg539_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg406_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg458_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg64_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg105_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg130_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add16_4_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_4_impl_0_out,
                 Y => Delay1No100_out);

SharedReg277_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg277_out;
SharedReg285_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg285_out;
SharedReg550_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg550_out;
SharedReg348_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg348_out;
SharedReg318_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg318_out;
SharedReg299_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg299_out;
SharedReg475_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg475_out;
SharedReg137_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg137_out;
SharedReg450_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg450_out;
SharedReg483_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg483_out;
SharedReg551_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg551_out;
SharedReg278_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg278_out;
SharedReg439_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg439_out;
SharedReg554_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg554_out;
SharedReg552_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg552_out;
SharedReg357_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg357_out;
   MUX_Add16_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg277_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg285_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg551_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg278_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg439_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg554_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg552_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg357_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg550_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg348_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg318_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg299_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg475_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg137_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg450_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg483_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add16_4_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_4_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Add17_4_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Add17_4_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Add17_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add17_4_impl_out,
                 X => Delay1No102_out_to_Add17_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Add17_4_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
SharedReg464_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg464_out;
SharedReg64_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg64_out;
SharedReg137_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg137_out;
SharedReg140_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg140_out;
SharedReg209_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg209_out;
SharedReg214_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg214_out;
SharedReg174_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg174_out;
Delay88No4_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_9_cast <= Delay88No4_out;
SharedReg540_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg540_out;
Delay111No4_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_11_cast <= Delay111No4_out;
   MUX_Add17_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg464_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay111No4_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg64_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg137_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg209_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg214_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg174_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay88No4_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg540_out_to_MUX_Add17_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add17_4_impl_0_LUT_out,
                 oMux => MUX_Add17_4_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add17_4_impl_0_out,
                 Y => Delay1No102_out);

SharedReg318_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg318_out;
SharedReg364_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg364_out;
SharedReg137_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg137_out;
SharedReg363_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg363_out;
SharedReg138_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg138_out;
SharedReg243_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg243_out;
SharedReg320_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg320_out;
SharedReg553_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg553_out;
Delay3No69_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_9_cast <= Delay3No69_out;
SharedReg372_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg372_out;
SharedReg535_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg535_out;
   MUX_Add17_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg318_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg364_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg535_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg137_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg363_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg138_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg243_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg320_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg553_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay3No69_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg372_out_to_MUX_Add17_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add17_4_impl_1_LUT_out,
                 oMux => MUX_Add17_4_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add17_4_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Add24_0_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Add24_0_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Add24_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add24_0_impl_out,
                 X => Delay1No104_out_to_Add24_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Add24_0_impl_parent_implementedSystem_port_1_cast);

SharedReg181_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg181_out;
SharedReg526_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg526_out;
Delay88No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_3_cast <= Delay88No_out;
SharedReg412_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg412_out;
Delay84No1_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_5_cast <= Delay84No1_out;
SharedReg36_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg36_out;
SharedReg19_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg19_out;
Delay43No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_8_cast <= Delay43No_out;
SharedReg413_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg413_out;
SharedReg47_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg47_out;
SharedReg533_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg533_out;
Delay90No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_12_cast <= Delay90No_out;
SharedReg411_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg411_out;
SharedReg507_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg507_out;
Delay41No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_15_cast <= Delay41No_out;
SharedReg89_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg89_out;
   MUX_Add24_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg181_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg526_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg533_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay90No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg411_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg507_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay41No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg89_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => Delay88No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg412_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay84No1_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg36_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg19_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay43No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg413_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg47_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add24_0_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add24_0_impl_0_out,
                 Y => Delay1No104_out);

SharedReg546_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg546_out;
SharedReg367_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg367_out;
SharedReg370_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg370_out;
SharedReg367_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg367_out;
SharedReg340_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg340_out;
SharedReg377_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg377_out;
SharedReg377_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg377_out;
SharedReg368_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg368_out;
SharedReg261_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg261_out;
SharedReg545_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg545_out;
SharedReg330_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg330_out;
SharedReg263_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg263_out;
SharedReg326_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg326_out;
SharedReg524_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg524_out;
SharedReg369_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg369_out;
SharedReg90_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg90_out;
   MUX_Add24_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg546_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg367_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg330_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg263_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg326_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg524_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg369_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg90_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg370_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg367_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg340_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg377_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg377_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg368_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg545_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Add24_0_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add24_0_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Add51_4_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Add51_4_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Add51_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add51_4_impl_out,
                 X => Delay1No106_out_to_Add51_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Add51_4_impl_parent_implementedSystem_port_1_cast);

SharedReg19_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg19_out;
SharedReg36_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg36_out;
SharedReg68_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg68_out;
Delay90No4_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_4_cast <= Delay90No4_out;
SharedReg448_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg448_out;
SharedReg447_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg447_out;
SharedReg515_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg515_out;
SharedReg468_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg468_out;
Delay32No4_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_9_cast <= Delay32No4_out;
Delay81No4_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_10_cast <= Delay81No4_out;
   MUX_Add51_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_10_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg19_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg36_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg68_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay90No4_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg448_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg447_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg515_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg468_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay32No4_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay81No4_out_to_MUX_Add51_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add51_4_impl_0_LUT_out,
                 oMux => MUX_Add51_4_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add51_4_impl_0_out,
                 Y => Delay1No106_out);

SharedReg553_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg553_out;
SharedReg361_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg361_out;
SharedReg376_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg376_out;
SharedReg353_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg353_out;
SharedReg319_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg319_out;
SharedReg372_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg372_out;
SharedReg374_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg374_out;
SharedReg551_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg551_out;
SharedReg535_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg535_out;
SharedReg541_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg541_out;
   MUX_Add51_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_10_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg553_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg361_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg376_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg319_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg372_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg374_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg551_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg535_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg541_out_to_MUX_Add51_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add51_4_impl_1_LUT_out,
                 oMux => MUX_Add51_4_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add51_4_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Product112_1_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Product112_1_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Product112_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product112_1_impl_out,
                 X => Delay1No108_out_to_Product112_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Product112_1_impl_parent_implementedSystem_port_1_cast);

SharedReg523_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg523_out;
SharedReg39_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg38_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg38_out;
SharedReg527_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg527_out;
SharedReg562_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg519_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg519_out;
SharedReg561_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg183_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg183_out;
SharedReg564_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg565_out;
SharedReg48_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg48_out;
SharedReg378_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg378_out;
SharedReg119_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg119_out;
SharedReg377_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg377_out;
SharedReg52_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg52_out;
   MUX_Product112_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg523_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg48_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg378_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg119_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg377_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg52_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg38_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg527_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg519_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg183_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product112_1_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_1_impl_0_out,
                 Y => Delay1No108_out);

SharedReg576_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg576_out;
SharedReg559_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg573_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg573_out;
SharedReg562_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg561_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg565_out;
SharedReg10_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg10_out;
SharedReg22_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg22_out;
SharedReg336_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg336_out;
SharedReg34_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg34_out;
SharedReg338_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg338_out;
   MUX_Product112_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg576_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg10_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg22_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg336_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg34_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg338_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg573_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product112_1_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_1_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Product112_2_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Product112_2_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Product112_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product112_2_impl_out,
                 X => Delay1No110_out_to_Product112_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Product112_2_impl_parent_implementedSystem_port_1_cast);

SharedReg54_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg54_out;
SharedReg504_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg504_out;
SharedReg499_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg499_out;
SharedReg294_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg294_out;
SharedReg37_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg37_out;
SharedReg31_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg31_out;
SharedReg385_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg385_out;
SharedReg562_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg499_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg499_out;
SharedReg561_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg156_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg156_out;
SharedReg564_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg565_out;
SharedReg76_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg76_out;
SharedReg386_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg386_out;
   MUX_Product112_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg54_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg504_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg156_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg564_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg565_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg76_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg386_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg499_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg294_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg37_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg31_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg385_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg499_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product112_2_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_2_impl_0_out,
                 Y => Delay1No110_out);

SharedReg33_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg33_out;
SharedReg578_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg578_out;
SharedReg570_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg570_out;
SharedReg347_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg347_out;
SharedReg559_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg14_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg14_out;
SharedReg573_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg573_out;
SharedReg562_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg563_out;
SharedReg561_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg565_out;
SharedReg10_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg10_out;
SharedReg22_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg22_out;
   MUX_Product112_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg33_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg578_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg564_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg565_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg10_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg22_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg570_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg347_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg14_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg573_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product112_2_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_2_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Product112_3_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Product112_3_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Product112_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product112_3_impl_out,
                 X => Delay1No112_out_to_Product112_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Product112_3_impl_parent_implementedSystem_port_1_cast);

SharedReg565_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg28_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg28_out;
SharedReg346_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg346_out;
SharedReg238_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg238_out;
SharedReg160_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg160_out;
SharedReg482_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg482_out;
SharedReg286_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg286_out;
SharedReg37_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg37_out;
SharedReg31_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg82_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg82_out;
SharedReg562_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg482_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg482_out;
SharedReg561_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg163_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg163_out;
SharedReg564_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg564_out;
   MUX_Product112_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg28_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg482_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg163_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg564_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg346_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg238_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg160_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg482_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg286_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg37_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg82_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product112_3_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_3_impl_0_out,
                 Y => Delay1No112_out);

SharedReg565_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg344_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg344_out;
SharedReg345_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg345_out;
SharedReg283_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg283_out;
SharedReg577_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg577_out;
SharedReg570_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg570_out;
SharedReg302_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg302_out;
SharedReg559_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg14_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg14_out;
SharedReg573_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg573_out;
SharedReg562_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg561_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg564_out;
   MUX_Product112_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg344_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg564_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg345_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg283_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg577_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg570_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg302_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg14_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg573_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product112_3_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_3_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Product113_4_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Product113_4_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Product113_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product113_4_impl_out,
                 X => Delay1No114_out_to_Product113_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Product113_4_impl_parent_implementedSystem_port_1_cast);

SharedReg561_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg131_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg131_out;
SharedReg458_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg458_out;
SharedReg564_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg299_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg299_out;
SharedReg393_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg393_out;
SharedReg238_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg238_out;
SharedReg130_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg130_out;
SharedReg458_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg458_out;
SharedReg402_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg402_out;
SharedReg7_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg7_out;
SharedReg400_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg400_out;
SharedReg561_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg236_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg236_out;
SharedReg236_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg236_out;
   MUX_Product113_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg131_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg7_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg400_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg236_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg236_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg458_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg299_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg393_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg238_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg130_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg458_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg402_out_to_MUX_Product113_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product113_4_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_4_impl_0_out,
                 Y => Delay1No114_out);

SharedReg561_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg566_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg566_out;
SharedReg564_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg28_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg28_out;
SharedReg29_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg29_out;
SharedReg22_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg22_out;
SharedReg569_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg569_out;
SharedReg570_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg570_out;
SharedReg374_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg374_out;
SharedReg13_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg13_out;
SharedReg572_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg572_out;
SharedReg561_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg564_out;
   MUX_Product113_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg13_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg572_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg564_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg566_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg28_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg29_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg22_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg569_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg570_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg374_out_to_MUX_Product113_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product113_4_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_4_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Product102_1_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Product102_1_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Product102_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product102_1_impl_out,
                 X => Delay1No116_out_to_Product102_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Product102_1_impl_parent_implementedSystem_port_1_cast);

Delay13No36_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_1_cast <= Delay13No36_out;
SharedReg7_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg7_out;
SharedReg425_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg425_out;
SharedReg561_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg215_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg215_out;
SharedReg215_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg215_out;
SharedReg565_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg176_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg176_out;
SharedReg519_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg519_out;
SharedReg367_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg367_out;
SharedReg12_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg12_out;
SharedReg18_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg18_out;
SharedReg219_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg219_out;
SharedReg180_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg180_out;
SharedReg507_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg507_out;
   MUX_Product102_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay13No36_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg367_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg12_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg18_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg219_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg180_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg507_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg425_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg215_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg215_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg176_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg519_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product102_1_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_1_impl_0_out,
                 Y => Delay1No116_out);

SharedReg576_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg576_out;
SharedReg13_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg572_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg572_out;
SharedReg561_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg16_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg16_out;
SharedReg566_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg566_out;
SharedReg17_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg17_out;
SharedReg367_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg367_out;
SharedReg369_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg369_out;
SharedReg576_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg576_out;
SharedReg578_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg578_out;
SharedReg570_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg570_out;
   MUX_Product102_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg576_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg17_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg367_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg369_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg576_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg578_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg570_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg572_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg16_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg566_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product102_1_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_1_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Product102_2_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Product102_2_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Product102_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product102_2_impl_out,
                 X => Delay1No118_out_to_Product102_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Product102_2_impl_parent_implementedSystem_port_1_cast);

SharedReg385_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg385_out;
SharedReg187_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg187_out;
SharedReg414_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg414_out;
SharedReg59_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg59_out;
SharedReg7_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg7_out;
SharedReg433_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg433_out;
SharedReg561_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg433_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg433_out;
SharedReg433_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg433_out;
SharedReg499_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg499_out;
SharedReg414_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg414_out;
SharedReg437_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg437_out;
SharedReg309_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg309_out;
SharedReg310_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg310_out;
SharedReg337_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg337_out;
   MUX_Product102_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg385_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg187_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg499_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg414_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg437_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg309_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg310_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg337_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg414_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg59_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg7_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg433_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg433_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg433_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product102_2_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_2_impl_0_out,
                 Y => Delay1No118_out);

SharedReg23_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg23_out;
SharedReg578_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg578_out;
SharedReg570_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg570_out;
SharedReg576_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg576_out;
SharedReg13_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg13_out;
SharedReg572_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg572_out;
SharedReg561_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg15_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg15_out;
SharedReg32_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg32_out;
SharedReg575_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg575_out;
SharedReg336_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg336_out;
SharedReg336_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg336_out;
SharedReg338_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg338_out;
   MUX_Product102_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg23_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg578_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg15_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg32_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg575_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg336_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg336_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg338_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg570_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg576_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg13_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg572_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product102_2_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_2_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Product102_3_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Product102_3_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Product102_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product102_3_impl_out,
                 X => Delay1No120_out_to_Product102_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Product102_3_impl_parent_implementedSystem_port_1_cast);

SharedReg565_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg12_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg12_out;
SharedReg18_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg18_out;
SharedReg107_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg107_out;
SharedReg99_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg99_out;
SharedReg419_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg419_out;
Delay13No38_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_7_cast <= Delay13No38_out;
SharedReg7_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg7_out;
SharedReg419_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg419_out;
SharedReg561_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg231_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg231_out;
SharedReg231_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg231_out;
SharedReg482_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg482_out;
SharedReg419_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg419_out;
SharedReg234_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg234_out;
   MUX_Product102_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg231_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg231_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg482_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg419_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg234_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg18_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg107_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg99_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg419_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay13No38_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg7_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg419_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product102_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product102_3_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_3_impl_0_out,
                 Y => Delay1No120_out);

SharedReg565_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg344_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg344_out;
SharedReg346_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg346_out;
SharedReg299_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg299_out;
SharedReg569_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg569_out;
SharedReg570_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg570_out;
SharedReg576_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg576_out;
SharedReg13_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg13_out;
SharedReg572_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg572_out;
SharedReg561_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg564_out;
SharedReg15_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg15_out;
SharedReg32_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg32_out;
SharedReg575_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg575_out;
   MUX_Product102_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg344_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg564_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg15_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg32_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg575_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg346_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg299_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg569_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg570_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg576_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg13_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg572_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product102_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product102_3_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_3_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Product104_0_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Product104_0_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Product104_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product104_0_impl_out,
                 X => Delay1No122_out_to_Product104_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Product104_0_impl_parent_implementedSystem_port_1_cast);

SharedReg527_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg527_out;
SharedReg1_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg141_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg141_out;
SharedReg175_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg175_out;
SharedReg565_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg508_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg508_out;
SharedReg407_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg407_out;
SharedReg507_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg507_out;
SharedReg367_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg367_out;
SharedReg176_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg176_out;
SharedReg329_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg329_out;
SharedReg407_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg407_out;
SharedReg407_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg407_out;
   MUX_Product104_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg527_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg507_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg367_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg176_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg329_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg407_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg407_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg8_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg141_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg175_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg508_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg407_out_to_MUX_Product104_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product104_0_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product104_0_impl_0_out,
                 Y => Delay1No122_out);

SharedReg571_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg571_out;
SharedReg20_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg27_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg27_out;
SharedReg566_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg566_out;
SharedReg567_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg567_out;
SharedReg28_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg28_out;
SharedReg29_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg29_out;
SharedReg24_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg24_out;
SharedReg569_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg569_out;
SharedReg570_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg570_out;
   MUX_Product104_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg571_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg567_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg28_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg29_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg24_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg569_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg570_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg26_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg27_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg566_out_to_MUX_Product104_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product104_0_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product104_0_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Product104_1_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Product104_1_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Product104_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product104_1_impl_out,
                 X => Delay1No124_out_to_Product104_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Product104_1_impl_parent_implementedSystem_port_1_cast);

SharedReg101_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg101_out;
SharedReg433_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg433_out;
SharedReg433_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg433_out;
SharedReg499_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg499_out;
SharedReg1_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg223_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg223_out;
SharedReg223_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg223_out;
SharedReg565_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg565_out;
SharedReg149_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg149_out;
SharedReg490_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg490_out;
SharedReg336_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg336_out;
SharedReg12_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg12_out;
SharedReg18_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg18_out;
   MUX_Product104_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg101_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg433_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg149_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg490_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg336_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg12_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg18_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg433_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg499_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg8_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg223_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg223_out_to_MUX_Product104_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product104_1_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product104_1_impl_0_out,
                 Y => Delay1No124_out);

SharedReg344_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg344_out;
SharedReg569_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg569_out;
SharedReg570_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg570_out;
SharedReg571_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg571_out;
SharedReg20_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg26_out;
SharedReg561_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg565_out;
SharedReg16_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg16_out;
SharedReg566_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg566_out;
SharedReg17_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg17_out;
SharedReg336_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg336_out;
SharedReg338_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg338_out;
   MUX_Product104_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg344_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg569_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg16_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg566_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg17_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg336_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg338_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg570_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg571_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg26_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product104_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product104_1_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product104_1_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Product104_4_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Product104_4_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Product104_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product104_4_impl_out,
                 X => Delay1No126_out_to_Product104_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Product104_4_impl_parent_implementedSystem_port_1_cast);

SharedReg535_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg535_out;
SharedReg562_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg169_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg169_out;
SharedReg516_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg516_out;
SharedReg565_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg565_out;
SharedReg138_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg138_out;
SharedReg541_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg541_out;
SharedReg536_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg536_out;
SharedReg513_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg513_out;
SharedReg374_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg374_out;
SharedReg362_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg362_out;
SharedReg541_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg541_out;
SharedReg513_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg513_out;
SharedReg439_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg439_out;
SharedReg1_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1_out;
SharedReg464_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg464_out;
   MUX_Product104_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg535_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg362_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg541_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg513_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg439_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg464_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg169_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg516_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg565_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg138_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg541_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg536_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg513_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg374_out_to_MUX_Product104_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product104_4_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product104_4_impl_0_out,
                 Y => Delay1No126_out);

SharedReg573_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg573_out;
SharedReg562_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg565_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg565_out;
SharedReg16_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg16_out;
SharedReg566_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg566_out;
SharedReg372_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg372_out;
SharedReg372_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg372_out;
SharedReg373_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg373_out;
SharedReg24_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg24_out;
SharedReg569_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg569_out;
SharedReg570_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg570_out;
SharedReg571_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg571_out;
SharedReg20_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg20_out;
SharedReg572_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg572_out;
   MUX_Product104_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg573_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg24_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg569_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg570_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg571_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg20_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg572_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg563_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg565_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg16_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg566_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg372_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg372_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg373_out_to_MUX_Product104_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product104_4_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product104_4_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Product105_2_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Product105_2_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Product105_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product105_2_impl_out,
                 X => Delay1No128_out_to_Product105_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Product105_2_impl_parent_implementedSystem_port_1_cast);

SharedReg565_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg292_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg292_out;
SharedReg345_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg345_out;
SharedReg392_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg392_out;
SharedReg196_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg196_out;
SharedReg449_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg449_out;
SharedReg286_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg286_out;
SharedReg25_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg25_out;
SharedReg482_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg482_out;
SharedReg561_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg419_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg419_out;
SharedReg482_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg482_out;
SharedReg234_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg234_out;
SharedReg449_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg449_out;
SharedReg482_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg482_out;
   MUX_Product105_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg292_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg419_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg482_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg234_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg449_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg482_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg345_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg392_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg196_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg449_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg286_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg25_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg482_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product105_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product105_2_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product105_2_impl_0_out,
                 Y => Delay1No128_out);

SharedReg565_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg344_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg344_out;
SharedReg346_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg346_out;
SharedReg23_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg23_out;
SharedReg578_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg578_out;
SharedReg570_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg570_out;
SharedReg35_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg35_out;
SharedReg20_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg20_out;
SharedReg572_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg572_out;
SharedReg561_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg564_out;
SharedReg574_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg574_out;
SharedReg3_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg3_out;
SharedReg566_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg566_out;
   MUX_Product105_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg344_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg564_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg574_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg3_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg566_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg346_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg23_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg578_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg570_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg35_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg20_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg572_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product105_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product105_2_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product105_2_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Product105_3_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Product105_3_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Product105_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product105_3_impl_out,
                 X => Delay1No130_out_to_Product105_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Product105_3_impl_parent_implementedSystem_port_1_cast);

SharedReg561_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg400_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg400_out;
SharedReg239_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg239_out;
SharedReg564_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg12_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg12_out;
SharedReg18_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg18_out;
SharedReg459_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg459_out;
SharedReg205_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg205_out;
SharedReg469_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg469_out;
SharedReg71_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg71_out;
SharedReg25_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg25_out;
SharedReg469_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg469_out;
SharedReg561_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg400_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg400_out;
SharedReg469_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg469_out;
   MUX_Product105_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg400_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg25_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg469_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg400_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg469_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg239_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg12_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg18_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg459_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg205_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg469_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg71_out_to_MUX_Product105_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product105_3_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product105_3_impl_0_out,
                 Y => Delay1No130_out);

SharedReg561_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg32_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg32_out;
SharedReg575_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg575_out;
SharedReg564_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg299_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg299_out;
SharedReg301_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg301_out;
SharedReg11_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg11_out;
SharedReg578_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg578_out;
SharedReg570_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg570_out;
SharedReg373_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg373_out;
SharedReg20_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg572_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg572_out;
SharedReg561_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg564_out;
   MUX_Product105_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg32_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg572_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg564_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg575_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg299_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg301_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg11_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg578_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg570_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg373_out_to_MUX_Product105_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product105_3_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product105_3_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Product105_4_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Product105_4_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Product105_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product105_4_impl_out,
                 X => Delay1No132_out_to_Product105_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Product105_4_impl_parent_implementedSystem_port_1_cast);

SharedReg7_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg7_out;
SharedReg170_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg170_out;
SharedReg516_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg516_out;
SharedReg209_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg209_out;
SharedReg513_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg513_out;
SharedReg243_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg243_out;
SharedReg516_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg516_out;
SharedReg362_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg362_out;
SharedReg372_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg372_out;
SharedReg562_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg562_out;
SharedReg565_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg565_out;
   MUX_Product105_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg7_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg170_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg565_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg516_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg209_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg513_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg243_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg516_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg362_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg372_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg562_out_to_MUX_Product105_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product105_4_impl_0_LUT_out,
                 oMux => MUX_Product105_4_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product105_4_impl_0_out,
                 Y => Delay1No132_out);

SharedReg13_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg13_out;
SharedReg24_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg27_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg27_out;
SharedReg28_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg28_out;
SharedReg569_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg569_out;
SharedReg563_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg570_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg570_out;
SharedReg562_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg565_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg565_out;
SharedReg567_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg567_out;
SharedReg572_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg572_out;
   MUX_Product105_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg13_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg572_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg27_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg28_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg569_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg570_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg565_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg567_out_to_MUX_Product105_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product105_4_impl_1_LUT_out,
                 oMux => MUX_Product105_4_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product105_4_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Product241_4_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Product241_4_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Product241_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product241_4_impl_out,
                 X => Delay1No134_out_to_Product241_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Product241_4_impl_parent_implementedSystem_port_1_cast);

SharedReg561_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg458_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg458_out;
SharedReg469_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg469_out;
SharedReg564_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg284_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg284_out;
SharedReg300_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg300_out;
SharedReg65_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg65_out;
SharedReg163_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg163_out;
SharedReg400_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg400_out;
SharedReg72_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg72_out;
SharedReg1_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg458_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg458_out;
SharedReg476_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg476_out;
   MUX_Product241_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg458_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg8_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg458_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg476_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg469_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg284_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg300_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg65_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg163_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg400_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg72_out_to_MUX_Product241_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product241_4_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product241_4_impl_0_out,
                 Y => Delay1No134_out);

SharedReg561_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg3_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg566_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg566_out;
SharedReg564_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg299_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg299_out;
SharedReg301_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg301_out;
SharedReg22_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg22_out;
SharedReg569_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg569_out;
SharedReg570_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg570_out;
SharedReg361_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg361_out;
SharedReg13_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg31_out;
SharedReg561_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg564_out;
   MUX_Product241_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg13_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg31_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg564_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg566_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg299_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg301_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg22_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg569_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg570_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg361_out_to_MUX_Product241_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product241_4_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product241_4_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Product321_4_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Product321_4_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Product321_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_4_impl_out,
                 X => Delay1No136_out_to_Product321_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Product321_4_impl_parent_implementedSystem_port_1_cast);

SharedReg561_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg476_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg476_out;
SharedReg476_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg476_out;
SharedReg70_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg70_out;
SharedReg12_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg12_out;
SharedReg285_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg285_out;
SharedReg169_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg169_out;
SharedReg165_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg165_out;
SharedReg476_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg476_out;
SharedReg459_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg459_out;
SharedReg37_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg37_out;
SharedReg31_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg31_out;
SharedReg70_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg70_out;
SharedReg562_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg469_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg469_out;
SharedReg560_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg560_out;
   MUX_Product321_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg476_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg37_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg31_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg70_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg469_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg560_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg476_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg70_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg12_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg285_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg169_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg165_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg476_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg459_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product321_4_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_4_impl_0_out,
                 Y => Delay1No136_out);

SharedReg561_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg3_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg566_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg566_out;
SharedReg564_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg299_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg299_out;
SharedReg300_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg300_out;
SharedReg11_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg11_out;
SharedReg577_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg577_out;
SharedReg570_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg570_out;
SharedReg373_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg373_out;
SharedReg559_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg14_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg14_out;
SharedReg573_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg573_out;
SharedReg562_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg560_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg560_out;
   MUX_Product321_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg14_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg573_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg560_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg566_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg299_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg300_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg11_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg577_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg570_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg373_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product321_4_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_4_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Product361_3_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Product361_3_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Product361_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product361_3_impl_out,
                 X => Delay1No138_out_to_Product361_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Product361_3_impl_parent_implementedSystem_port_1_cast);

SharedReg83_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg83_out;
SharedReg12_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg12_out;
SharedReg293_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg293_out;
SharedReg201_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg201_out;
SharedReg123_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg123_out;
SharedReg231_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg231_out;
SharedReg6_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg6_out;
SharedReg1_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg449_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg449_out;
SharedReg392_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg392_out;
SharedReg395_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg395_out;
SharedReg392_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg392_out;
SharedReg392_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg392_out;
   MUX_Product361_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg83_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg449_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg392_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg395_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg392_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg392_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg293_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg201_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg123_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg231_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg6_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg8_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product361_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product361_3_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product361_3_impl_0_out,
                 Y => Delay1No138_out);

SharedReg9_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg344_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg344_out;
SharedReg345_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg345_out;
SharedReg299_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg299_out;
SharedReg569_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg569_out;
SharedReg570_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg570_out;
SharedReg302_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg302_out;
SharedReg13_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg561_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg564_out;
SharedReg574_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg574_out;
SharedReg3_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg3_out;
SharedReg566_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg566_out;
   MUX_Product361_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg344_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg564_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg574_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg3_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg566_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg345_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg299_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg569_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg570_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg302_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg13_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product361_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product361_3_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product361_3_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Product391_2_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Product391_2_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Product391_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product391_2_impl_out,
                 X => Delay1No140_out_to_Product391_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Product391_2_impl_parent_implementedSystem_port_1_cast);

SharedReg192_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg192_out;
SharedReg414_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg414_out;
SharedReg223_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg223_out;
SharedReg294_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg294_out;
SharedReg25_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg25_out;
SharedReg490_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg490_out;
SharedReg561_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg414_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg414_out;
SharedReg499_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg499_out;
SharedReg225_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg225_out;
SharedReg490_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg490_out;
SharedReg499_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg499_out;
SharedReg433_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg433_out;
SharedReg12_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg12_out;
SharedReg311_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg311_out;
   MUX_Product391_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg192_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg414_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg225_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg490_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg499_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg433_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg12_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg311_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg223_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg294_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg25_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg490_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg414_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg499_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product391_2_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product391_2_impl_0_out,
                 Y => Delay1No140_out);

SharedReg344_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg344_out;
SharedReg569_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg569_out;
SharedReg570_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg570_out;
SharedReg35_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg35_out;
SharedReg20_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg572_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg572_out;
SharedReg561_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg574_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg574_out;
SharedReg3_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg3_out;
SharedReg566_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg566_out;
SharedReg567_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg567_out;
SharedReg336_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg336_out;
SharedReg337_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg337_out;
   MUX_Product391_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg344_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg569_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg574_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg3_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg566_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg567_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg336_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg337_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg570_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg35_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg572_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product391_2_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product391_2_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Product441_2_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Product441_2_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Product441_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product441_2_impl_out,
                 X => Delay1No142_out_to_Product441_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Product441_2_impl_parent_implementedSystem_port_1_cast);

SharedReg233_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg233_out;
SharedReg153_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg153_out;
SharedReg490_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg490_out;
SharedReg6_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg6_out;
SharedReg1_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg490_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg490_out;
SharedReg385_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg385_out;
SharedReg502_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg502_out;
SharedReg385_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg385_out;
SharedReg385_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg385_out;
SharedReg4_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg4_out;
SharedReg28_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg28_out;
SharedReg338_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg338_out;
   MUX_Product441_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg233_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg153_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg502_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg385_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg385_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg4_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg28_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg338_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg490_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg6_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg8_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg490_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg385_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product441_2_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product441_2_impl_0_out,
                 Y => Delay1No142_out);

SharedReg291_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg291_out;
SharedReg577_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg577_out;
SharedReg570_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg570_out;
SharedReg347_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg347_out;
SharedReg13_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg31_out;
SharedReg561_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg574_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg574_out;
SharedReg3_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg3_out;
SharedReg566_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg566_out;
SharedReg336_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg336_out;
SharedReg336_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg336_out;
SharedReg337_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg337_out;
   MUX_Product441_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg291_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg577_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg574_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg3_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg566_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg336_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg336_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg337_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg570_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg347_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg13_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg31_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product441_2_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product441_2_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Product491_0_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Product491_0_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Product491_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product491_0_impl_out,
                 X => Delay1No144_out_to_Product491_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Product491_0_impl_parent_implementedSystem_port_1_cast);

SharedReg312_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg312_out;
SharedReg25_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg25_out;
SharedReg507_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg507_out;
SharedReg561_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg425_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg425_out;
SharedReg425_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg425_out;
SharedReg527_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg527_out;
SharedReg507_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg507_out;
SharedReg427_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg427_out;
SharedReg326_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg326_out;
SharedReg327_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg327_out;
SharedReg368_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg368_out;
SharedReg329_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg329_out;
SharedReg507_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg507_out;
SharedReg425_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg425_out;
   MUX_Product491_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg312_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg25_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg326_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg327_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg368_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg329_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg507_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg425_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg507_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg425_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg425_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg527_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg507_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg427_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product491_0_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product491_0_impl_0_out,
                 Y => Delay1No144_out);

SharedReg35_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg35_out;
SharedReg20_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg572_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg572_out;
SharedReg561_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg15_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg15_out;
SharedReg32_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg32_out;
SharedReg575_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg575_out;
SharedReg367_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg367_out;
SharedReg367_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg367_out;
SharedReg369_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg369_out;
SharedReg35_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg35_out;
SharedReg569_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg569_out;
SharedReg570_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg570_out;
   MUX_Product491_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg35_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg367_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg367_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg369_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg35_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg569_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg570_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg572_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg15_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg32_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg575_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product491_0_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product491_0_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Product512_4_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Product512_4_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Product512_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product512_4_impl_out,
                 X => Delay1No146_out_to_Product512_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Product512_4_impl_parent_implementedSystem_port_1_cast);

SharedReg12_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg12_out;
SharedReg8_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
SharedReg25_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg25_out;
SharedReg477_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg477_out;
SharedReg464_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg464_out;
SharedReg248_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg248_out;
SharedReg246_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg246_out;
SharedReg439_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg439_out;
SharedReg372_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg372_out;
SharedReg565_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg565_out;
SharedReg562_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
   MUX_Product512_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg12_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg25_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg477_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg464_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg248_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg246_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg439_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg372_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg565_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product512_4_impl_0_LUT_out,
                 oMux => MUX_Product512_4_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_4_impl_0_out,
                 Y => Delay1No146_out);

SharedReg16_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg16_out;
SharedReg17_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg20_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg31_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg31_out;
SharedReg372_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg372_out;
SharedReg562_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg562_out;
SharedReg565_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg565_out;
SharedReg570_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg570_out;
SharedReg578_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg578_out;
SharedReg576_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg576_out;
SharedReg563_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg563_out;
   MUX_Product512_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg16_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg563_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg20_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg31_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg372_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg562_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg565_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg570_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg578_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg576_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product512_4_impl_1_LUT_out,
                 oMux => MUX_Product512_4_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_4_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Product55_4_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Product55_4_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Product55_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_4_impl_out,
                 X => Delay1No148_out_to_Product55_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Product55_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg31_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg31_out;
SharedReg513_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg513_out;
SharedReg243_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg243_out;
SharedReg535_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg535_out;
SharedReg516_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg516_out;
SharedReg464_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg464_out;
SharedReg360_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg360_out;
SharedReg362_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg362_out;
SharedReg359_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg359_out;
SharedReg562_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
   MUX_Product55_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg513_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg243_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg535_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg516_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg464_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg360_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg362_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg359_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product55_4_impl_0_LUT_out,
                 oMux => MUX_Product55_4_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_4_impl_0_out,
                 Y => Delay1No148_out);

SharedReg15_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg14_out;
SharedReg13_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg13_out;
SharedReg32_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg32_out;
SharedReg35_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg35_out;
SharedReg372_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg372_out;
SharedReg372_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg372_out;
SharedReg562_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg570_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg570_out;
SharedReg569_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg569_out;
SharedReg563_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg563_out;
   MUX_Product55_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg15_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg14_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg563_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg13_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg32_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg35_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg372_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg372_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg570_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg569_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product55_4_impl_1_LUT_out,
                 oMux => MUX_Product55_4_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_4_impl_1_out,
                 Y => Delay1No149_out);

Delay1No150_out_to_Product56_0_impl_parent_implementedSystem_port_0_cast <= Delay1No150_out;
Delay1No151_out_to_Product56_0_impl_parent_implementedSystem_port_1_cast <= Delay1No151_out;
   Product56_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product56_0_impl_out,
                 X => Delay1No150_out_to_Product56_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No151_out_to_Product56_0_impl_parent_implementedSystem_port_1_cast);

SharedReg6_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg6_out;
SharedReg1_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg407_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg407_out;
SharedReg519_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg519_out;
SharedReg218_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg218_out;
SharedReg519_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg519_out;
SharedReg527_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg527_out;
SharedReg407_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg407_out;
SharedReg12_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg12_out;
SharedReg328_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg328_out;
SharedReg520_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg520_out;
SharedReg511_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg511_out;
SharedReg519_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg519_out;
   MUX_Product56_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg6_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg407_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg12_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg328_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg520_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg511_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg519_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg8_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg407_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg519_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg218_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg519_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg527_out_to_MUX_Product56_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product56_0_impl_0_out);

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product56_0_impl_0_out,
                 Y => Delay1No150_out);

SharedReg339_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg339_out;
SharedReg13_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg31_out;
SharedReg561_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg574_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg574_out;
SharedReg3_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg3_out;
SharedReg566_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg566_out;
SharedReg567_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg567_out;
SharedReg367_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg367_out;
SharedReg368_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg368_out;
SharedReg568_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg568_out;
SharedReg577_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg577_out;
SharedReg570_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg570_out;
   MUX_Product56_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg339_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg567_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg367_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg368_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg568_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg577_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg570_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg31_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg574_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg3_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg566_out_to_MUX_Product56_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product56_0_impl_1_out);

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product56_0_impl_1_out,
                 Y => Delay1No151_out);

Delay1No152_out_to_Product611_0_impl_parent_implementedSystem_port_0_cast <= Delay1No152_out;
Delay1No153_out_to_Product611_0_impl_parent_implementedSystem_port_1_cast <= Delay1No153_out;
   Product611_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product611_0_impl_out,
                 X => Delay1No152_out_to_Product611_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No153_out_to_Product611_0_impl_parent_implementedSystem_port_1_cast);

SharedReg312_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg312_out;
SharedReg37_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg37_out;
SharedReg31_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg31_out;
SharedReg561_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg507_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg507_out;
SharedReg527_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg527_out;
SharedReg521_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg521_out;
SharedReg377_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg377_out;
SharedReg377_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg377_out;
SharedReg4_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg4_out;
SharedReg28_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg28_out;
SharedReg369_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg369_out;
SharedReg529_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg529_out;
SharedReg523_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg523_out;
SharedReg527_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg527_out;
   MUX_Product611_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg312_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg37_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg4_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg28_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg369_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg529_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg523_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg527_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg31_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg507_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg527_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg521_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg377_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg377_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product611_0_impl_0_out);

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product611_0_impl_0_out,
                 Y => Delay1No152_out);

SharedReg339_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg339_out;
SharedReg559_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg14_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg14_out;
SharedReg561_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg563_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg574_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg574_out;
SharedReg3_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg3_out;
SharedReg566_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg566_out;
SharedReg367_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg367_out;
SharedReg367_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg367_out;
SharedReg368_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg368_out;
SharedReg568_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg568_out;
SharedReg578_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg578_out;
SharedReg570_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg570_out;
   MUX_Product611_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg339_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg367_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg367_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg368_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg568_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg578_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg570_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg14_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg574_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg3_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg566_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Product611_0_impl_1_out);

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product611_0_impl_1_out,
                 Y => Delay1No153_out);

Delay1No154_out_to_Product611_4_impl_parent_implementedSystem_port_0_cast <= Delay1No154_out;
Delay1No155_out_to_Product611_4_impl_parent_implementedSystem_port_1_cast <= Delay1No155_out;
   Product611_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product611_4_impl_out,
                 X => Delay1No154_out_to_Product611_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No155_out_to_Product611_4_impl_parent_implementedSystem_port_1_cast);

SharedReg12_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg12_out;
SharedReg37_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg37_out;
SharedReg38_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg38_out;
SharedReg516_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg516_out;
SharedReg443_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg443_out;
SharedReg541_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg541_out;
Delay14No24_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_7_cast <= Delay14No24_out;
SharedReg169_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg169_out;
SharedReg245_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg245_out;
SharedReg513_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg513_out;
SharedReg562_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
   MUX_Product611_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg12_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg37_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg38_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg516_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg443_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg541_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay14No24_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg169_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg245_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg513_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product611_4_impl_0_LUT_out,
                 oMux => MUX_Product611_4_impl_0_out);

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product611_4_impl_0_out,
                 Y => Delay1No154_out);

SharedReg3_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg3_out;
SharedReg372_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg372_out;
SharedReg568_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg568_out;
SharedReg559_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg559_out;
SharedReg570_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg562_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg562_out;
SharedReg574_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg574_out;
SharedReg567_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg567_out;
SharedReg577_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg577_out;
SharedReg560_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg560_out;
   MUX_Product611_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg3_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg372_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg560_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg568_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg559_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg570_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg562_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg574_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg567_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg577_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product611_4_impl_1_LUT_out,
                 oMux => MUX_Product611_4_impl_1_out);

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product611_4_impl_1_out,
                 Y => Delay1No155_out);

Delay1No156_out_to_Product811_4_impl_parent_implementedSystem_port_0_cast <= Delay1No156_out;
Delay1No157_out_to_Product811_4_impl_parent_implementedSystem_port_1_cast <= Delay1No157_out;
   Product811_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product811_4_impl_out,
                 X => Delay1No156_out_to_Product811_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No157_out_to_Product811_4_impl_parent_implementedSystem_port_1_cast);

SharedReg4_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg4_out;
SharedReg28_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg28_out;
SharedReg39_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg39_out;
SharedReg541_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg541_out;
SharedReg517_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg517_out;
SharedReg538_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg538_out;
SharedReg442_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg442_out;
SharedReg516_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg516_out;
SharedReg562_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg562_out;
   MUX_Product811_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg4_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg28_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg39_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg541_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg517_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg538_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg442_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg516_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg562_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_Product811_4_impl_0_LUT_out,
                 oMux => MUX_Product811_4_impl_0_out);

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product811_4_impl_0_out,
                 Y => Delay1No156_out);

SharedReg3_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg3_out;
SharedReg372_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg372_out;
SharedReg372_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg372_out;
SharedReg568_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg568_out;
SharedReg578_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg578_out;
SharedReg563_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg562_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg562_out;
SharedReg574_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg574_out;
SharedReg559_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg559_out;
   MUX_Product811_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg3_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg372_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg372_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg568_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg578_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg562_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg574_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg559_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_9_cast,
                 iSel => MUX_Product811_4_impl_1_LUT_out,
                 oMux => MUX_Product811_4_impl_1_out);

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product811_4_impl_1_out,
                 Y => Delay1No157_out);

Delay1No158_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No158_out;
Delay1No159_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No159_out;
   Subtract12_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_0_impl_out,
                 X => Delay1No158_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No159_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg129_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg129_out;
SharedReg43_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg43_out;
SharedReg115_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg115_out;
SharedReg428_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg428_out;
SharedReg92_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg92_out;
SharedReg116_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg116_out;
SharedReg46_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg46_out;
SharedReg510_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg510_out;
SharedReg116_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg116_out;
SharedReg179_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg179_out;
Delay33No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_11_cast <= Delay33No_out;
SharedReg429_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg429_out;
SharedReg432_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg432_out;
Delay33No1_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_14_cast <= Delay33No1_out;
SharedReg222_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg222_out;
SharedReg230_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg230_out;
   MUX_Subtract12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg129_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg43_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay33No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg429_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg432_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay33No1_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg222_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg230_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg115_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg428_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg92_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg116_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg46_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg510_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg116_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg179_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Subtract12_0_impl_0_out);

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_0_impl_0_out,
                 Y => Delay1No158_out);

SharedReg270_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg270_out;
SharedReg326_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg326_out;
SharedReg251_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg251_out;
SharedReg252_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg252_out;
SharedReg367_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg367_out;
SharedReg251_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg251_out;
SharedReg328_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg328_out;
SharedReg253_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg253_out;
SharedReg262_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg262_out;
SharedReg330_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg330_out;
SharedReg253_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg253_out;
SharedReg329_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg329_out;
SharedReg371_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg371_out;
SharedReg262_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg262_out;
SharedReg251_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg251_out;
SharedReg340_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg340_out;
   MUX_Subtract12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg270_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg326_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg253_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg329_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg371_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg262_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg251_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg340_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg251_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg252_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg367_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg251_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg328_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg253_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg262_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg330_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Subtract12_0_impl_1_out);

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_0_impl_1_out,
                 Y => Delay1No159_out);

Delay1No160_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No160_out;
Delay1No161_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No161_out;
   Subtract12_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_1_impl_out,
                 X => Delay1No160_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No161_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg134_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg134_out;
SharedReg189_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg189_out;
Delay64No2_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast <= Delay64No2_out;
SharedReg136_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg136_out;
SharedReg379_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg379_out;
SharedReg97_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg97_out;
SharedReg226_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg226_out;
SharedReg51_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg51_out;
SharedReg98_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg98_out;
SharedReg381_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg381_out;
SharedReg417_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg417_out;
SharedReg98_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg98_out;
SharedReg152_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg152_out;
SharedReg424_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg424_out;
SharedReg438_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg438_out;
SharedReg388_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg388_out;
   MUX_Subtract12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg134_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg189_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg417_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg98_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg152_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg424_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg438_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg388_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => Delay64No2_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg136_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg379_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg97_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg226_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg51_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg98_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg381_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Subtract12_1_impl_0_out);

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_1_impl_0_out,
                 Y => Delay1No160_out);

SharedReg286_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg286_out;
SharedReg259_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg259_out;
SharedReg348_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg348_out;
SharedReg279_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg279_out;
SharedReg309_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg309_out;
SharedReg309_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg309_out;
SharedReg261_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg261_out;
SharedReg268_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg268_out;
SharedReg259_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg259_out;
SharedReg338_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg338_out;
SharedReg312_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg312_out;
SharedReg270_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg270_out;
SharedReg313_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg313_out;
SharedReg294_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg294_out;
SharedReg312_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg312_out;
SharedReg295_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg295_out;
   MUX_Subtract12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg286_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg259_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg312_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg270_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg313_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg294_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg312_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg295_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg348_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg279_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg309_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg309_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg261_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg268_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg259_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg338_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Subtract12_1_impl_1_out);

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_1_impl_1_out,
                 Y => Delay1No161_out);

Delay1No162_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No162_out;
Delay1No163_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No163_out;
   Subtract12_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_2_impl_out,
                 X => Delay1No162_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No163_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast);

SharedReg466_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg466_out;
SharedReg423_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg423_out;
SharedReg86_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg86_out;
SharedReg403_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg403_out;
SharedReg161_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg161_out;
Delay64No3_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_6_cast <= Delay64No3_out;
SharedReg247_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg247_out;
SharedReg436_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg436_out;
SharedReg57_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg57_out;
SharedReg193_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg193_out;
SharedReg56_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg56_out;
SharedReg58_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg58_out;
SharedReg80_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg80_out;
SharedReg108_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg108_out;
SharedReg102_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg102_out;
SharedReg62_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg62_out;
   MUX_Subtract12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg466_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg423_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg56_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg58_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg80_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg108_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg102_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg62_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg86_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg403_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg161_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay64No3_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg247_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg436_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg57_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg193_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Subtract12_2_impl_0_out);

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_2_impl_0_out,
                 Y => Delay1No162_out);

SharedReg319_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg319_out;
SharedReg294_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg294_out;
SharedReg287_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg287_out;
SharedReg319_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg319_out;
SharedReg268_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg268_out;
SharedReg303_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg303_out;
SharedReg303_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg303_out;
SharedReg344_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg344_out;
SharedReg291_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg291_out;
SharedReg293_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg293_out;
SharedReg276_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg276_out;
SharedReg268_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg268_out;
SharedReg346_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg346_out;
SharedReg353_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg353_out;
SharedReg279_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg279_out;
SharedReg301_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg301_out;
   MUX_Subtract12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_16_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg319_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg294_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg276_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg268_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg346_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg353_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg279_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg301_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_2 => SharedReg287_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg319_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg268_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg303_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg303_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg344_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg291_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg293_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount161_out,
                 oMux => MUX_Subtract12_2_impl_1_out);

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_2_impl_1_out,
                 Y => Delay1No163_out);

Delay1No164_out_to_Subtract12_3_impl_parent_implementedSystem_port_0_cast <= Delay1No164_out;
Delay1No165_out_to_Subtract12_3_impl_parent_implementedSystem_port_1_cast <= Delay1No165_out;
   Subtract12_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_3_impl_out,
                 X => Delay1No164_out_to_Subtract12_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No165_out_to_Subtract12_3_impl_parent_implementedSystem_port_1_cast);

SharedReg404_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg404_out;
SharedReg444_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg444_out;
SharedReg421_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg421_out;
SharedReg110_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg110_out;
SharedReg172_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg172_out;
SharedReg133_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg133_out;
SharedReg172_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg172_out;
SharedReg109_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg109_out;
SharedReg474_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg474_out;
SharedReg240_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg240_out;
SharedReg167_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg167_out;
Delay64No4_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_12_cast <= Delay64No4_out;
   MUX_Subtract12_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg404_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg444_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg167_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay64No4_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg421_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg110_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg172_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg133_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg172_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg109_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg474_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg240_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Subtract12_3_impl_0_LUT_out,
                 oMux => MUX_Subtract12_3_impl_0_out);

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_3_impl_0_out,
                 Y => Delay1No164_out);

SharedReg276_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg276_out;
SharedReg283_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg283_out;
SharedReg283_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg283_out;
SharedReg299_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg299_out;
SharedReg285_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg285_out;
SharedReg283_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg283_out;
SharedReg286_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg286_out;
SharedReg362_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg362_out;
SharedReg299_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg299_out;
SharedReg355_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg355_out;
SharedReg320_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg320_out;
SharedReg376_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg376_out;
   MUX_Subtract12_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg276_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg283_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg320_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg376_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg283_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg299_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg285_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg283_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg286_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg362_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg299_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg355_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Subtract12_3_impl_1_LUT_out,
                 oMux => MUX_Subtract12_3_impl_1_out);

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_3_impl_1_out,
                 Y => Delay1No165_out);

Delay1No166_out_to_Subtract10_4_impl_parent_implementedSystem_port_0_cast <= Delay1No166_out;
Delay1No167_out_to_Subtract10_4_impl_parent_implementedSystem_port_1_cast <= Delay1No167_out;
   Subtract10_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract10_4_impl_out,
                 X => Delay1No166_out_to_Subtract10_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No167_out_to_Subtract10_4_impl_parent_implementedSystem_port_1_cast);

SharedReg461_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg461_out;
SharedReg66_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg518_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg518_out;
Delay22No4_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_4_cast <= Delay22No4_out;
SharedReg75_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg75_out;
   MUX_Subtract10_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg461_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg518_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay22No4_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg75_out_to_MUX_Subtract10_4_impl_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Subtract10_4_impl_0_LUT_out,
                 oMux => MUX_Subtract10_4_impl_0_out);

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_4_impl_0_out,
                 Y => Delay1No166_out);

SharedReg355_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg355_out;
SharedReg318_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg318_out;
SharedReg355_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg355_out;
SharedReg359_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg359_out;
SharedReg359_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg359_out;
   MUX_Subtract10_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg355_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg318_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg355_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg359_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg359_out_to_MUX_Subtract10_4_impl_1_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Subtract10_4_impl_1_LUT_out,
                 oMux => MUX_Subtract10_4_impl_1_out);

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_4_impl_1_out,
                 Y => Delay1No167_out);
   Constant1_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);

Delay1No168_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast <= Delay1No168_out;
Delay1No169_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast <= Delay1No169_out;
   Divide_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Divide_0_impl_out,
                 X => Delay1No168_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No169_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast);

SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg555_out;
SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg555_out;
SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg555_out;
SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg555_out;
SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg555_out;
   MUX_Divide_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg555_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Divide_0_impl_0_LUT_out,
                 oMux => MUX_Divide_0_impl_0_out);

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Divide_0_impl_0_out,
                 Y => Delay1No168_out);

SharedReg367_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg367_out;
SharedReg336_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg336_out;
SharedReg276_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg276_out;
SharedReg283_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg283_out;
SharedReg372_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg372_out;
   MUX_Divide_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg367_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg336_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg276_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg283_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg372_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Divide_0_impl_1_LUT_out,
                 oMux => MUX_Divide_0_impl_1_out);

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Divide_0_impl_1_out,
                 Y => Delay1No169_out);
   Constant_0_impl_instance: Constant_float_8_23_348_mult_8en9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);

   Delay133No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => Delay133No_out);

   Delay133No1_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => Delay133No1_out);

   Delay133No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => Delay133No2_out);

   Delay133No4_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => Delay133No4_out);

   Delay131No4_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => Delay131No4_out);

   Delay125No3_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => Delay125No3_out);

   Delay130No_instance: Delay_34_DelayLength_125_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=125 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg371_out,
                 Y => Delay130No_out);

   Delay130No1_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => Delay130No1_out);

   Delay130No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => Delay130No2_out);

   Delay130No3_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => Delay130No3_out);

   Delay130No4_instance: Delay_34_DelayLength_125_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=125 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => Delay130No4_out);

   Delay133No5_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg335_out,
                 Y => Delay133No5_out);

   Delay133No6_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => Delay133No6_out);

   Delay133No7_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => Delay133No7_out);

   Delay133No9_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => Delay133No9_out);

   Delay25No_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => Delay25No_out);

   Delay11No40_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => Delay11No40_out);

   Delay19No2_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => Delay19No2_out);

   Delay19No4_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => Delay19No4_out);

   Delay21No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => Delay21No_out);

   Delay22No4_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => Delay22No4_out);

   Delay13No30_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => Delay13No30_out);

   Delay16No17_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => Delay16No17_out);

   Delay33No_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => Delay33No_out);

   Delay33No1_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => Delay33No1_out);

   Delay13No36_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => Delay13No36_out);

   Delay13No38_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => Delay13No38_out);

   Delay2No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg550_out,
                 Y => Delay2No132_out);

   Delay3No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg546_out,
                 Y => Delay3No65_out);

   Delay3No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg554_out,
                 Y => Delay3No69_out);

   Delay14No16_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => Delay14No16_out);

   Delay88No_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg526_out,
                 Y => Delay88No_out);

   Delay88No1_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg498_out,
                 Y => Delay88No1_out);

   Delay88No3_instance: Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=63 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => Delay88No3_out);

   Delay88No4_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg540_out,
                 Y => Delay88No4_out);

   Delay80No3_instance: Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=37 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => Delay80No3_out);

   Delay84No_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg432_out,
                 Y => Delay84No_out);

   Delay84No1_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => Delay84No1_out);

   Delay84No2_instance: Delay_34_DelayLength_71_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=71 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => Delay84No2_out);

   Delay84No3_instance: Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=68 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => Delay84No3_out);

   Delay84No4_instance: Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=43 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg468_out,
                 Y => Delay84No4_out);

   Delay90No_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg413_out,
                 Y => Delay90No_out);

   Delay90No1_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => Delay90No1_out);

   Delay90No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg457_out,
                 Y => Delay90No2_out);

   Delay90No3_instance: Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=49 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg463_out,
                 Y => Delay90No3_out);

   Delay90No4_instance: Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=55 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg515_out,
                 Y => Delay90No4_out);

   Delay67No2_instance: Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=54 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg424_out,
                 Y => Delay67No2_out);

   Delay67No3_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg406_out,
                 Y => Delay67No3_out);

   Delay59No_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => Delay59No_out);

   Delay59No2_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => Delay59No2_out);

   Delay64No2_instance: Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=41 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => Delay64No2_out);

   Delay64No3_instance: Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=46 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => Delay64No3_out);

   Delay64No4_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => Delay64No4_out);

   Delay35No1_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => Delay35No1_out);

   Delay35No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => Delay35No2_out);

   Delay35No3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => Delay35No3_out);

   Delay14No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg518_out,
                 Y => Delay14No24_out);

   Delay41No_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg512_out,
                 Y => Delay41No_out);

   Delay43No_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => Delay43No_out);

   Delay43No1_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => Delay43No1_out);

   Delay43No2_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => Delay43No2_out);

   Delay43No4_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => Delay43No4_out);

   Delay32No1_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg438_out,
                 Y => Delay32No1_out);

   Delay32No2_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => Delay32No2_out);

   Delay32No4_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => Delay32No4_out);

   Delay81No1_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg391_out,
                 Y => Delay81No1_out);

   Delay81No2_instance: Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=65 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => Delay81No2_out);

   Delay81No3_instance: Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=48 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => Delay81No3_out);

   Delay81No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg544_out,
                 Y => Delay81No4_out);

   Delay111No_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg534_out,
                 Y => Delay111No_out);

   Delay111No1_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg506_out,
                 Y => Delay111No1_out);

   Delay111No2_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg489_out,
                 Y => Delay111No2_out);

   Delay111No3_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg481_out,
                 Y => Delay111No3_out);

   Delay111No4_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg448_out,
                 Y => Delay111No4_out);

   MUX_Inv_11_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Inv_11_0_0_LUT_out);

   MUX_Inv_12_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Inv_12_0_0_LUT_out);

   MUX_Inv_13_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Inv_13_0_0_LUT_out);

   MUX_Inv_21_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Inv_21_0_0_LUT_out);

   MUX_Inv_22_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Inv_22_0_0_LUT_out);

   MUX_Inv_23_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Inv_23_0_0_LUT_out);

   MUX_Inv_31_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Inv_31_0_0_LUT_out);

   MUX_Inv_32_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Inv_32_0_0_LUT_out);

   MUX_Inv_33_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Inv_33_0_0_LUT_out);

   MUX_Inv_41_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Inv_41_0_0_LUT_out);

   MUX_Inv_42_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Inv_42_0_0_LUT_out);

   MUX_Inv_43_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Inv_43_0_0_LUT_out);

   MUX_Add17_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add17_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Add17_4_impl_0_LUT_out);

   MUX_Add17_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add17_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Add17_4_impl_1_LUT_out);

   MUX_Add51_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add51_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Add51_4_impl_0_LUT_out);

   MUX_Add51_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add51_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Add51_4_impl_1_LUT_out);

   MUX_Product105_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product105_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Product105_4_impl_0_LUT_out);

   MUX_Product105_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product105_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Product105_4_impl_1_LUT_out);

   MUX_Product512_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product512_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Product512_4_impl_0_LUT_out);

   MUX_Product512_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product512_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Product512_4_impl_1_LUT_out);

   MUX_Product55_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product55_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Product55_4_impl_0_LUT_out);

   MUX_Product55_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product55_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Product55_4_impl_1_LUT_out);

   MUX_Product611_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product611_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Product611_4_impl_0_LUT_out);

   MUX_Product611_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product611_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Product611_4_impl_1_LUT_out);

   MUX_Product811_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Product811_4_impl_0_LUT_out);

   MUX_Product811_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Product811_4_impl_1_LUT_out);

   MUX_Subtract12_3_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract12_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Subtract12_3_impl_0_LUT_out);

   MUX_Subtract12_3_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract12_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Subtract12_3_impl_1_LUT_out);

   MUX_Subtract10_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract10_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Subtract10_4_impl_0_LUT_out);

   MUX_Subtract10_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract10_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Subtract10_4_impl_1_LUT_out);

   MUX_Divide_0_impl_0_LUT_instance: GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Divide_0_impl_0_LUT_out);

   MUX_Divide_0_impl_1_LUT_instance: GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount161_out,
                 Output => MUX_Divide_0_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_0_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg2_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg3_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg4_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_0_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg7_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg8_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg9_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg10_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg11_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_0_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg13_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg14_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg15_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg16_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg17_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_0_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_0_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg20_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg21_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg22_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg23_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_0_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg25_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg26_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg27_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg28_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_0_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg30_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg31_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_0_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_0_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_0_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_0_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_0_impl_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_1_impl_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_2_impl_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_3_impl_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_4_impl_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_4_impl_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_2_impl_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_3_impl_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_0_impl_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_1_impl_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_2_impl_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_3_impl_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_0_impl_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_1_impl_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_2_impl_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_3_impl_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_4_impl_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_0_impl_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_1_impl_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_2_impl_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_3_impl_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_4_impl_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_0_impl_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_1_impl_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_2_impl_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_3_impl_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_4_impl_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_0_impl_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_1_impl_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=46 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_2_impl_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_3_impl_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_4_impl_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_0_impl_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=99 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_1_impl_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_98_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=98 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg263_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_2_impl_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_98_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=98 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_3_impl_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_98_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=98 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_4_impl_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_123_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=123 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_2_impl_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_108_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=108 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_4_impl_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_94_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=94 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add101_1_impl_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_94_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=94 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_4_impl_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_98_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=98 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add141_0_impl_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_94_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=94 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg332_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg334_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add151_2_impl_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_119_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=119 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg341_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add151_3_impl_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg344_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg346_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=104 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg349_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add16_4_impl_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg353_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=107 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg357_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add17_4_impl_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg359_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg360_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg361_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg362_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_108_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=108 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg365_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add24_0_impl_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg368_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg369_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add51_4_impl_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg372_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg375_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product112_1_impl_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg377_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg380_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product112_2_impl_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg385_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg387_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg388_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg389_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg390_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product112_3_impl_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg396_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product113_4_impl_out,
                 Y => SharedReg400_out);

   SharedReg401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => SharedReg401_out);

   SharedReg402_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg401_out,
                 Y => SharedReg402_out);

   SharedReg403_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg402_out,
                 Y => SharedReg403_out);

   SharedReg404_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg403_out,
                 Y => SharedReg404_out);

   SharedReg405_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg404_out,
                 Y => SharedReg405_out);

   SharedReg406_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg405_out,
                 Y => SharedReg406_out);

   SharedReg407_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product102_1_impl_out,
                 Y => SharedReg407_out);

   SharedReg408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg407_out,
                 Y => SharedReg408_out);

   SharedReg409_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => SharedReg409_out);

   SharedReg410_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg409_out,
                 Y => SharedReg410_out);

   SharedReg411_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg410_out,
                 Y => SharedReg411_out);

   SharedReg412_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg411_out,
                 Y => SharedReg412_out);

   SharedReg413_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg412_out,
                 Y => SharedReg413_out);

   SharedReg414_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product102_2_impl_out,
                 Y => SharedReg414_out);

   SharedReg415_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg414_out,
                 Y => SharedReg415_out);

   SharedReg416_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg415_out,
                 Y => SharedReg416_out);

   SharedReg417_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg416_out,
                 Y => SharedReg417_out);

   SharedReg418_instance: Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=54 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg417_out,
                 Y => SharedReg418_out);

   SharedReg419_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product102_3_impl_out,
                 Y => SharedReg419_out);

   SharedReg420_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg419_out,
                 Y => SharedReg420_out);

   SharedReg421_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => SharedReg421_out);

   SharedReg422_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg421_out,
                 Y => SharedReg422_out);

   SharedReg423_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg422_out,
                 Y => SharedReg423_out);

   SharedReg424_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg423_out,
                 Y => SharedReg424_out);

   SharedReg425_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product104_0_impl_out,
                 Y => SharedReg425_out);

   SharedReg426_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg425_out,
                 Y => SharedReg426_out);

   SharedReg427_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg426_out,
                 Y => SharedReg427_out);

   SharedReg428_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg427_out,
                 Y => SharedReg428_out);

   SharedReg429_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => SharedReg429_out);

   SharedReg430_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg429_out,
                 Y => SharedReg430_out);

   SharedReg431_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg430_out,
                 Y => SharedReg431_out);

   SharedReg432_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg431_out,
                 Y => SharedReg432_out);

   SharedReg433_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product104_1_impl_out,
                 Y => SharedReg433_out);

   SharedReg434_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg433_out,
                 Y => SharedReg434_out);

   SharedReg435_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg434_out,
                 Y => SharedReg435_out);

   SharedReg436_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg435_out,
                 Y => SharedReg436_out);

   SharedReg437_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg436_out,
                 Y => SharedReg437_out);

   SharedReg438_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg437_out,
                 Y => SharedReg438_out);

   SharedReg439_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product104_4_impl_out,
                 Y => SharedReg439_out);

   SharedReg440_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => SharedReg440_out);

   SharedReg441_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg440_out,
                 Y => SharedReg441_out);

   SharedReg442_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg441_out,
                 Y => SharedReg442_out);

   SharedReg443_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => SharedReg443_out);

   SharedReg444_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg443_out,
                 Y => SharedReg444_out);

   SharedReg445_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg444_out,
                 Y => SharedReg445_out);

   SharedReg446_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg445_out,
                 Y => SharedReg446_out);

   SharedReg447_instance: Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=46 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg446_out,
                 Y => SharedReg447_out);

   SharedReg448_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg447_out,
                 Y => SharedReg448_out);

   SharedReg449_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product105_2_impl_out,
                 Y => SharedReg449_out);

   SharedReg450_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg449_out,
                 Y => SharedReg450_out);

   SharedReg451_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg450_out,
                 Y => SharedReg451_out);

   SharedReg452_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg451_out,
                 Y => SharedReg452_out);

   SharedReg453_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg452_out,
                 Y => SharedReg453_out);

   SharedReg454_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg453_out,
                 Y => SharedReg454_out);

   SharedReg455_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg454_out,
                 Y => SharedReg455_out);

   SharedReg456_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg455_out,
                 Y => SharedReg456_out);

   SharedReg457_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg456_out,
                 Y => SharedReg457_out);

   SharedReg458_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product105_3_impl_out,
                 Y => SharedReg458_out);

   SharedReg459_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg458_out,
                 Y => SharedReg459_out);

   SharedReg460_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg459_out,
                 Y => SharedReg460_out);

   SharedReg461_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg460_out,
                 Y => SharedReg461_out);

   SharedReg462_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg461_out,
                 Y => SharedReg462_out);

   SharedReg463_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg462_out,
                 Y => SharedReg463_out);

   SharedReg464_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product105_4_impl_out,
                 Y => SharedReg464_out);

   SharedReg465_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg464_out,
                 Y => SharedReg465_out);

   SharedReg466_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg465_out,
                 Y => SharedReg466_out);

   SharedReg467_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg466_out,
                 Y => SharedReg467_out);

   SharedReg468_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg467_out,
                 Y => SharedReg468_out);

   SharedReg469_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product241_4_impl_out,
                 Y => SharedReg469_out);

   SharedReg470_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg469_out,
                 Y => SharedReg470_out);

   SharedReg471_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg470_out,
                 Y => SharedReg471_out);

   SharedReg472_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg471_out,
                 Y => SharedReg472_out);

   SharedReg473_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg472_out,
                 Y => SharedReg473_out);

   SharedReg474_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg473_out,
                 Y => SharedReg474_out);

   SharedReg475_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg474_out,
                 Y => SharedReg475_out);

   SharedReg476_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_4_impl_out,
                 Y => SharedReg476_out);

   SharedReg477_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg476_out,
                 Y => SharedReg477_out);

   SharedReg478_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg477_out,
                 Y => SharedReg478_out);

   SharedReg479_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg478_out,
                 Y => SharedReg479_out);

   SharedReg480_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg479_out,
                 Y => SharedReg480_out);

   SharedReg481_instance: Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=43 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg480_out,
                 Y => SharedReg481_out);

   SharedReg482_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product361_3_impl_out,
                 Y => SharedReg482_out);

   SharedReg483_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg482_out,
                 Y => SharedReg483_out);

   SharedReg484_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg483_out,
                 Y => SharedReg484_out);

   SharedReg485_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg484_out,
                 Y => SharedReg485_out);

   SharedReg486_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg485_out,
                 Y => SharedReg486_out);

   SharedReg487_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg486_out,
                 Y => SharedReg487_out);

   SharedReg488_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg487_out,
                 Y => SharedReg488_out);

   SharedReg489_instance: Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=61 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg488_out,
                 Y => SharedReg489_out);

   SharedReg490_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product391_2_impl_out,
                 Y => SharedReg490_out);

   SharedReg491_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg490_out,
                 Y => SharedReg491_out);

   SharedReg492_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg491_out,
                 Y => SharedReg492_out);

   SharedReg493_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg492_out,
                 Y => SharedReg493_out);

   SharedReg494_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg493_out,
                 Y => SharedReg494_out);

   SharedReg495_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg494_out,
                 Y => SharedReg495_out);

   SharedReg496_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg495_out,
                 Y => SharedReg496_out);

   SharedReg497_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg496_out,
                 Y => SharedReg497_out);

   SharedReg498_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg497_out,
                 Y => SharedReg498_out);

   SharedReg499_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product441_2_impl_out,
                 Y => SharedReg499_out);

   SharedReg500_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg499_out,
                 Y => SharedReg500_out);

   SharedReg501_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg500_out,
                 Y => SharedReg501_out);

   SharedReg502_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg501_out,
                 Y => SharedReg502_out);

   SharedReg503_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg502_out,
                 Y => SharedReg503_out);

   SharedReg504_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg503_out,
                 Y => SharedReg504_out);

   SharedReg505_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg504_out,
                 Y => SharedReg505_out);

   SharedReg506_instance: Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=64 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg505_out,
                 Y => SharedReg506_out);

   SharedReg507_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product491_0_impl_out,
                 Y => SharedReg507_out);

   SharedReg508_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg507_out,
                 Y => SharedReg508_out);

   SharedReg509_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg508_out,
                 Y => SharedReg509_out);

   SharedReg510_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg509_out,
                 Y => SharedReg510_out);

   SharedReg511_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg510_out,
                 Y => SharedReg511_out);

   SharedReg512_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg511_out,
                 Y => SharedReg512_out);

   SharedReg513_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product512_4_impl_out,
                 Y => SharedReg513_out);

   SharedReg514_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg513_out,
                 Y => SharedReg514_out);

   SharedReg515_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg514_out,
                 Y => SharedReg515_out);

   SharedReg516_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_4_impl_out,
                 Y => SharedReg516_out);

   SharedReg517_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg516_out,
                 Y => SharedReg517_out);

   SharedReg518_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg517_out,
                 Y => SharedReg518_out);

   SharedReg519_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product56_0_impl_out,
                 Y => SharedReg519_out);

   SharedReg520_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg519_out,
                 Y => SharedReg520_out);

   SharedReg521_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg520_out,
                 Y => SharedReg521_out);

   SharedReg522_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg521_out,
                 Y => SharedReg522_out);

   SharedReg523_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg522_out,
                 Y => SharedReg523_out);

   SharedReg524_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg523_out,
                 Y => SharedReg524_out);

   SharedReg525_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg524_out,
                 Y => SharedReg525_out);

   SharedReg526_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg525_out,
                 Y => SharedReg526_out);

   SharedReg527_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product611_0_impl_out,
                 Y => SharedReg527_out);

   SharedReg528_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg527_out,
                 Y => SharedReg528_out);

   SharedReg529_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg528_out,
                 Y => SharedReg529_out);

   SharedReg530_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg529_out,
                 Y => SharedReg530_out);

   SharedReg531_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg530_out,
                 Y => SharedReg531_out);

   SharedReg532_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => SharedReg532_out);

   SharedReg533_instance: Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=62 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg532_out,
                 Y => SharedReg533_out);

   SharedReg534_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg533_out,
                 Y => SharedReg534_out);

   SharedReg535_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product611_4_impl_out,
                 Y => SharedReg535_out);

   SharedReg536_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg535_out,
                 Y => SharedReg536_out);

   SharedReg537_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg536_out,
                 Y => SharedReg537_out);

   SharedReg538_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg537_out,
                 Y => SharedReg538_out);

   SharedReg539_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg538_out,
                 Y => SharedReg539_out);

   SharedReg540_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg539_out,
                 Y => SharedReg540_out);

   SharedReg541_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product811_4_impl_out,
                 Y => SharedReg541_out);

   SharedReg542_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg541_out,
                 Y => SharedReg542_out);

   SharedReg543_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg542_out,
                 Y => SharedReg543_out);

   SharedReg544_instance: Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=62 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg543_out,
                 Y => SharedReg544_out);

   SharedReg545_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_0_impl_out,
                 Y => SharedReg545_out);

   SharedReg546_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg545_out,
                 Y => SharedReg546_out);

   SharedReg547_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_1_impl_out,
                 Y => SharedReg547_out);

   SharedReg548_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg547_out,
                 Y => SharedReg548_out);

   SharedReg549_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg548_out,
                 Y => SharedReg549_out);

   SharedReg550_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_2_impl_out,
                 Y => SharedReg550_out);

   SharedReg551_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_3_impl_out,
                 Y => SharedReg551_out);

   SharedReg552_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg551_out,
                 Y => SharedReg552_out);

   SharedReg553_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract10_4_impl_out,
                 Y => SharedReg553_out);

   SharedReg554_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg553_out,
                 Y => SharedReg554_out);

   SharedReg555_instance: Delay_34_DelayLength_144_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=144 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg555_out);

   SharedReg556_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Divide_0_impl_out,
                 Y => SharedReg556_out);

   SharedReg557_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg556_out,
                 Y => SharedReg557_out);

   SharedReg558_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg557_out,
                 Y => SharedReg558_out);

   SharedReg559_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg559_out);

   SharedReg560_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg559_out,
                 Y => SharedReg560_out);

   SharedReg561_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg560_out,
                 Y => SharedReg561_out);

   SharedReg562_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg561_out,
                 Y => SharedReg562_out);

   SharedReg563_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg562_out,
                 Y => SharedReg563_out);

   SharedReg564_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg563_out,
                 Y => SharedReg564_out);

   SharedReg565_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg564_out,
                 Y => SharedReg565_out);

   SharedReg566_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg565_out,
                 Y => SharedReg566_out);

   SharedReg567_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg566_out,
                 Y => SharedReg567_out);

   SharedReg568_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg567_out,
                 Y => SharedReg568_out);

   SharedReg569_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg568_out,
                 Y => SharedReg569_out);

   SharedReg570_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg569_out,
                 Y => SharedReg570_out);

   SharedReg571_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg570_out,
                 Y => SharedReg571_out);

   SharedReg572_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg571_out,
                 Y => SharedReg572_out);

   SharedReg573_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg572_out,
                 Y => SharedReg573_out);

   SharedReg574_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg573_out,
                 Y => SharedReg574_out);

   SharedReg575_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg574_out,
                 Y => SharedReg575_out);

   SharedReg576_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg575_out,
                 Y => SharedReg576_out);

   SharedReg577_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg576_out,
                 Y => SharedReg577_out);

   SharedReg578_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg577_out,
                 Y => SharedReg578_out);
end architecture;

