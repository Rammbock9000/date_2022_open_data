--------------------------------------------------------------------------------
--                         ModuloCounter_64_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_64_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of ModuloCounter_64_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(5 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 63 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1942393
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1942393 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1942393 is
signal XX_m1942394 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m1942394 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m1942394 <= X ;
   YY_m1942394 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid1942397
--                   (IntAdderClassical_33_f500_uid1942399)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid1942397 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid1942397 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1942393 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid1942397 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1942393  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
   RoundingAdder: IntAdder_33_f500_uid1942397  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound   ,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_64_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_64_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iS_51 : in std_logic_vector(33 downto 0);
          iS_52 : in std_logic_vector(33 downto 0);
          iS_53 : in std_logic_vector(33 downto 0);
          iS_54 : in std_logic_vector(33 downto 0);
          iS_55 : in std_logic_vector(33 downto 0);
          iS_56 : in std_logic_vector(33 downto 0);
          iS_57 : in std_logic_vector(33 downto 0);
          iS_58 : in std_logic_vector(33 downto 0);
          iS_59 : in std_logic_vector(33 downto 0);
          iS_60 : in std_logic_vector(33 downto 0);
          iS_61 : in std_logic_vector(33 downto 0);
          iS_62 : in std_logic_vector(33 downto 0);
          iS_63 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_64_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
         iS_51 when "110011",
         iS_52 when "110100",
         iS_53 when "110101",
         iS_54 when "110110",
         iS_55 when "110111",
         iS_56 when "111000",
         iS_57 when "111001",
         iS_58 when "111010",
         iS_59 when "111011",
         iS_60 when "111100",
         iS_61 when "111101",
         iS_62 when "111110",
         iS_63 when "111111",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid1942458_RightShifter
--                (RightShifter_24_by_max_26_F250_uid1942460)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1942458_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1942458_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid1942463
--                  (IntAdderAlternative_27_f250_uid1942467)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid1942463 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid1942463 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid1942470
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid1942470 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid1942470 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid1942473
--                   (IntAdderClassical_34_f250_uid1942475)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid1942473 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid1942473 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid1942458
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1942458 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1942458 is
   component FPAdd_8_23_uid1942458_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid1942463 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid1942470 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid1942473 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid1942458_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid1942463  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid1942470  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid1942473  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid1942458 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid1942458  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_61_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_61_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iS_51 : in std_logic_vector(33 downto 0);
          iS_52 : in std_logic_vector(33 downto 0);
          iS_53 : in std_logic_vector(33 downto 0);
          iS_54 : in std_logic_vector(33 downto 0);
          iS_55 : in std_logic_vector(33 downto 0);
          iS_56 : in std_logic_vector(33 downto 0);
          iS_57 : in std_logic_vector(33 downto 0);
          iS_58 : in std_logic_vector(33 downto 0);
          iS_59 : in std_logic_vector(33 downto 0);
          iS_60 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_61_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
         iS_51 when "110011",
         iS_52 when "110100",
         iS_53 when "110101",
         iS_54 when "110110",
         iS_55 when "110111",
         iS_56 when "111000",
         iS_57 when "111001",
         iS_58 when "111010",
         iS_59 when "111011",
         iS_60 when "111100",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_34_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_34_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_34_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_51_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_51_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_51_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_20_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_20_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(4 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_20_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00000",
         iS_1 when "00001",
         iS_2 when "00010",
         iS_3 when "00011",
         iS_4 when "00100",
         iS_5 when "00101",
         iS_6 when "00110",
         iS_7 when "00111",
         iS_8 when "01000",
         iS_9 when "01001",
         iS_10 when "01010",
         iS_11 when "01011",
         iS_12 when "01100",
         iS_13 when "01101",
         iS_14 when "01110",
         iS_15 when "01111",
         iS_16 when "10000",
         iS_17 when "10001",
         iS_18 when "10010",
         iS_19 when "10011",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_13_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_13_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_13_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
         iS_11 when "1011",
         iS_12 when "1100",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_6_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_6_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_6_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
         iS_5 when "101",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_3_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_3_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(1 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_3_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00",
         iS_1 when "01",
         iS_2 when "10",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_2_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(0 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0",
         iS_1 when "1",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_0_617123672897668340553423149685841053724_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_617123672897668340553423149685841053724_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_617123672897668340553423149685841053724_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111000111011111101111010001";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_0_631862801488796588245122620719484984875_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_631862801488796588245122620719484984875_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_631862801488796588245122620719484984875_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001000011100000111000011";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_1_436934552725145586293820088030770421028_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_436934552725145586293820088030770421028_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_436934552725145586293820088030770421028_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111101101111110110101111001";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_1_561088850170149200380365073215216398239_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_561088850170149200380365073215216398239_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_561088850170149200380365073215216398239_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111110001111101000111000010";
end architecture;

--------------------------------------------------------------------------------
--   Constant_float_8_23_1_67381401040949318037576176720904186368_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_67381401040949318037576176720904186368_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_67381401040949318037576176720904186368_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111110101100011111110001010";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_1_767419732788928943278961014584638178349_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_767419732788928943278961014584638178349_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_767419732788928943278961014584638178349_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111111000100011101011001111";
end architecture;

--------------------------------------------------------------------------------
--   Constant_float_8_23_1_83466961525726479642628419242100790143_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_83466961525726479642628419242100790143_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_83466961525726479642628419242100790143_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111111010101101011001110100";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_1_869869533302351394254969818575773388147_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_869869533302351394254969818575773388147_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_869869533302351394254969818575773388147_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111111011110101011111100011";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_0_663686724095854829741369940165895968676_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_663686724095854829741369940165895968676_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_663686724095854829741369940165895968676_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001010011110011101100000";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_0_712333225863809871292176012502750381827_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_712333225863809871292176012502750381827_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_712333225863809871292176012502750381827_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001101100101101101111000";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_0_777424256340159325340266605053329840302_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_777424256340159325340266605053329840302_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_777424256340159325340266605053329840302_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111010001110000010101000111";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_0_858338451424324633265428019512910395861_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_858338451424324633265428019512910395861_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_858338451424324633265428019512910395861_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111010110111011110000010010";
end architecture;

--------------------------------------------------------------------------------
--   Constant_float_8_23_0_95403875322976861017565397560247220099_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_95403875322976861017565397560247220099_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_95403875322976861017565397560247220099_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111011101000011101111100010";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_1_062858000783881262663044253713451325893_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_062858000783881262663044253713451325893_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_062858000783881262663044253713451325893_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100010000000101110111011";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_1_182256984960216694702239692560397088528_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_182256984960216694702239692560397088528_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_182256984960216694702239692560397088528_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100101110101010000110010";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_1_308589307952890523623068474989850074053_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_308589307952890523623068474989850074053_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_308589307952890523623068474989850074053_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111101001110111111111011011";
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0101000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_99584180311675085661704542872030287981_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_99584180311675085661704542872030287981_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_99584180311675085661704542872030287981_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011111101110111101111101";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_987534845729581944873132215434452518821_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_987534845729581944873132215434452518821_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_987534845729581944873132215434452518821_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011111001100111100010101";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_906979034015293006376623452524654567242_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_906979034015293006376623452524654567242_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_906979034015293006376623452524654567242_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011010000010111111000111";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_898568629504465254953515795932617038488_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_898568629504465254953515795932617038488_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_898568629504465254953515795932617038488_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011001100000100010011000";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_891139475905879052675118145998567342758_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_891139475905879052675118145998567342758_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_891139475905879052675118145998567342758_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011001000010000110110111";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_885091234632599865861379839770961552858_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_885091234632599865861379839770961552858_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_885091234632599865861379839770961552858_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011000101001010101010111";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_880803415623673480183697392931208014488_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_880803415623673480183697392931208014488_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_880803415623673480183697392931208014488_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011000010111110001010101";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_878576235602384070233483726042322814465_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_878576235602384070233483726042322814465_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_878576235602384070233483726042322814465_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011000001110101001011111";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_979173278459382512295405831537209451199_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_979173278459382512295405831537209451199_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_979173278459382512295405831537209451199_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011110101010101100011010";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_970685163049390786760284299816703423858_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_970685163049390786760284299816703423858_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_970685163049390786760284299816703423858_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011110000111111011010011";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_962013487567665803723571116279345005751_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_962013487567665803723571116279345005751_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_962013487567665803723571116279345005751_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011101100100011010000100";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_95312319664069156122110371143207885325_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_95312319664069156122110371143207885325_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_95312319664069156122110371143207885325_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011100111111111111100010";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_944010225685960935315677033941028639674_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_944010225685960935315677033941028639674_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_944010225685960935315677033941028639674_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011100011010101010100111";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_934712586109242460352675152535084635019_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_934712586109242460352675152535084635019_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_934712586109242460352675152535084635019_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011110100100101010011";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_925322845902050161726037913467735052109_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_925322845902050161726037913467735052109_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_925322845902050161726037913467735052109_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001110000111110101";
end architecture;

--------------------------------------------------------------------------------
--  Constant_float_8_23_n0_916000226493365876656582713621901348233_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n0_916000226493365876656582713621901348233_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n0_916000226493365876656582713621901348233_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011010100111111011111110";
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 37 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      Y <= s36;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 22 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      Y <= s21;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum1_0_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum1_0_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum1_0_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "110111" when "000000",
      "000000" when "000001",
      "011100" when "000010",
      "110101" when "000011",
      "000000" when "000100",
      "010010" when "000101",
      "011111" when "000110",
      "001010" when "000111",
      "101101" when "001000",
      "011110" when "001001",
      "010000" when "001010",
      "010110" when "001011",
      "100101" when "001100",
      "000111" when "001101",
      "000101" when "001110",
      "000010" when "001111",
      "001000" when "010000",
      "100111" when "010001",
      "100011" when "010010",
      "100001" when "010011",
      "111011" when "010100",
      "101000" when "010101",
      "000000" when "010110",
      "010011" when "010111",
      "001110" when "011000",
      "101010" when "011001",
      "010001" when "011010",
      "011000" when "011011",
      "001011" when "011100",
      "101100" when "011101",
      "011010" when "011110",
      "111001" when "011111",
      "010101" when "100000",
      "101111" when "100001",
      "010111" when "100010",
      "110010" when "100011",
      "000011" when "100100",
      "110100" when "100101",
      "000000" when "100110",
      "110110" when "100111",
      "100010" when "101000",
      "111100" when "101001",
      "101001" when "101010",
      "111000" when "101011",
      "010100" when "101100",
      "011101" when "101101",
      "101011" when "101110",
      "000100" when "101111",
      "011001" when "110000",
      "100000" when "110001",
      "111010" when "110010",
      "011011" when "110011",
      "110001" when "110100",
      "001111" when "110101",
      "110000" when "110110",
      "001100" when "110111",
      "110011" when "111000",
      "000110" when "111001",
      "101110" when "111010",
      "001001" when "111011",
      "100110" when "111100",
      "100100" when "111101",
      "000001" when "111110",
      "001101" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum1_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum1_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum1_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Sum1_0_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum1_0_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum1_0_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum1_0_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum1_0_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "111001" when "000000",
      "000000" when "000001",
      "011100" when "000010",
      "110000" when "000011",
      "000000" when "000100",
      "010010" when "000101",
      "100000" when "000110",
      "001001" when "000111",
      "101100" when "001000",
      "011111" when "001001",
      "010000" when "001010",
      "010110" when "001011",
      "101000" when "001100",
      "001100" when "001101",
      "000101" when "001110",
      "000010" when "001111",
      "000111" when "010000",
      "101010" when "010001",
      "110010" when "010010",
      "100100" when "010011",
      "100010" when "010100",
      "100110" when "010101",
      "000000" when "010110",
      "010011" when "010111",
      "001110" when "011000",
      "111011" when "011001",
      "010001" when "011010",
      "011000" when "011011",
      "001010" when "011100",
      "101011" when "011101",
      "011010" when "011110",
      "101110" when "011111",
      "010101" when "100000",
      "110100" when "100001",
      "010111" when "100010",
      "110110" when "100011",
      "000011" when "100100",
      "101111" when "100101",
      "000000" when "100110",
      "110001" when "100111",
      "100101" when "101000",
      "100011" when "101001",
      "100111" when "101010",
      "111010" when "101011",
      "010100" when "101100",
      "011101" when "101101",
      "111100" when "101110",
      "000100" when "101111",
      "011001" when "110000",
      "100001" when "110001",
      "011110" when "110010",
      "011011" when "110011",
      "111000" when "110100",
      "001111" when "110101",
      "110101" when "110110",
      "001011" when "110111",
      "110111" when "111000",
      "000110" when "111001",
      "101101" when "111010",
      "001000" when "111011",
      "101001" when "111100",
      "110011" when "111101",
      "000001" when "111110",
      "001101" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum1_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum1_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum1_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Sum1_0_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum1_0_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum1_1_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum1_1_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum1_1_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000000" when "000000",
      "000000" when "000001",
      "001100" when "000010",
      "000000" when "000011",
      "000000" when "000100",
      "000000" when "000101",
      "000000" when "000110",
      "100001" when "000111",
      "000000" when "001000",
      "011100" when "001001",
      "100000" when "001010",
      "000000" when "001011",
      "010100" when "001100",
      "000000" when "001101",
      "011101" when "001110",
      "000000" when "001111",
      "000000" when "010000",
      "011001" when "010001",
      "011110" when "010010",
      "000001" when "010011",
      "001000" when "010100",
      "000000" when "010101",
      "000000" when "010110",
      "010010" when "010111",
      "010101" when "011000",
      "011010" when "011001",
      "010000" when "011010",
      "000000" when "011011",
      "000000" when "011100",
      "000000" when "011101",
      "000111" when "011110",
      "010110" when "011111",
      "001010" when "100000",
      "000000" when "100001",
      "000110" when "100010",
      "010111" when "100011",
      "000000" when "100100",
      "011011" when "100101",
      "000000" when "100110",
      "001110" when "100111",
      "000000" when "101000",
      "000010" when "101001",
      "000100" when "101010",
      "000000" when "101011",
      "000000" when "101100",
      "010011" when "101101",
      "000000" when "101110",
      "001011" when "101111",
      "000000" when "110000",
      "000000" when "110001",
      "000101" when "110010",
      "000000" when "110011",
      "011111" when "110100",
      "001101" when "110101",
      "000000" when "110110",
      "001001" when "110111",
      "000000" when "111000",
      "000000" when "111001",
      "000011" when "111010",
      "000000" when "111011",
      "011000" when "111100",
      "000000" when "111101",
      "001111" when "111110",
      "010001" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum1_1_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum1_1_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum1_1_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Sum1_1_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum1_1_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum1_1_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum1_1_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum1_1_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000000" when "000000",
      "000000" when "000001",
      "001100" when "000010",
      "000000" when "000011",
      "011000" when "000100",
      "000000" when "000101",
      "000000" when "000110",
      "010101" when "000111",
      "000000" when "001000",
      "100001" when "001001",
      "011100" when "001010",
      "000000" when "001011",
      "010001" when "001100",
      "000000" when "001101",
      "100000" when "001110",
      "000000" when "001111",
      "000000" when "010000",
      "011111" when "010001",
      "011101" when "010010",
      "000000" when "010011",
      "000111" when "010100",
      "000000" when "010101",
      "000000" when "010110",
      "010010" when "010111",
      "010100" when "011000",
      "010110" when "011001",
      "001011" when "011010",
      "000000" when "011011",
      "000000" when "011100",
      "000000" when "011101",
      "000110" when "011110",
      "010111" when "011111",
      "001001" when "100000",
      "000000" when "100001",
      "000101" when "100010",
      "011001" when "100011",
      "000000" when "100100",
      "011010" when "100101",
      "000000" when "100110",
      "001111" when "100111",
      "000000" when "101000",
      "000001" when "101001",
      "000011" when "101010",
      "000000" when "101011",
      "000000" when "101100",
      "010011" when "101101",
      "000000" when "101110",
      "001010" when "101111",
      "000000" when "110000",
      "000000" when "110001",
      "000100" when "110010",
      "000000" when "110011",
      "011011" when "110100",
      "001101" when "110101",
      "000000" when "110110",
      "001000" when "110111",
      "000000" when "111000",
      "000000" when "111001",
      "000010" when "111010",
      "000000" when "111011",
      "011110" when "111100",
      "000000" when "111101",
      "001110" when "111110",
      "010000" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum1_1_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum1_1_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum1_1_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Sum1_1_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum1_1_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum1_2_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum1_2_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum1_2_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "100011" when "000000",
      "000000" when "000001",
      "011000" when "000010",
      "001101" when "000011",
      "100010" when "000100",
      "000000" when "000101",
      "010001" when "000110",
      "011001" when "000111",
      "000000" when "001000",
      "001010" when "001001",
      "010100" when "001010",
      "101110" when "001011",
      "001001" when "001100",
      "010000" when "001101",
      "011110" when "001110",
      "100101" when "001111",
      "101000" when "010000",
      "110001" when "010001",
      "001110" when "010010",
      "000010" when "010011",
      "010101" when "010100",
      "101111" when "010101",
      "000000" when "010110",
      "101001" when "010111",
      "101011" when "011000",
      "000001" when "011001",
      "000011" when "011010",
      "011100" when "011011",
      "011010" when "011100",
      "110010" when "011101",
      "011011" when "011110",
      "100110" when "011111",
      "101101" when "100000",
      "100001" when "100001",
      "000101" when "100010",
      "000100" when "100011",
      "000000" when "100100",
      "001000" when "100101",
      "000000" when "100110",
      "100000" when "100111",
      "000000" when "101000",
      "010110" when "101001",
      "001011" when "101010",
      "000000" when "101011",
      "101010" when "101100",
      "001100" when "101101",
      "101100" when "101110",
      "010010" when "101111",
      "000000" when "110000",
      "000000" when "110001",
      "100100" when "110010",
      "000000" when "110011",
      "011101" when "110100",
      "010011" when "110101",
      "000000" when "110110",
      "010111" when "110111",
      "000110" when "111000",
      "011111" when "111001",
      "100111" when "111010",
      "000000" when "111011",
      "110000" when "111100",
      "001111" when "111101",
      "000000" when "111110",
      "000111" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum1_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum1_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum1_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Sum1_2_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum1_2_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum1_2_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum1_2_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum1_2_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "011101" when "000000",
      "000000" when "000001",
      "011000" when "000010",
      "001101" when "000011",
      "011100" when "000100",
      "000000" when "000101",
      "010000" when "000110",
      "110001" when "000111",
      "000000" when "001000",
      "001000" when "001001",
      "010100" when "001010",
      "101100" when "001011",
      "000111" when "001100",
      "001111" when "001101",
      "100000" when "001110",
      "100110" when "001111",
      "101000" when "010000",
      "100100" when "010001",
      "010010" when "010010",
      "000010" when "010011",
      "010101" when "010100",
      "110000" when "010101",
      "000000" when "010110",
      "101110" when "010111",
      "101001" when "011000",
      "000001" when "011001",
      "000011" when "011010",
      "011011" when "011011",
      "110010" when "011100",
      "011001" when "011101",
      "011010" when "011110",
      "101101" when "011111",
      "100010" when "100000",
      "011111" when "100001",
      "001001" when "100010",
      "000100" when "100011",
      "000000" when "100100",
      "000110" when "100101",
      "000000" when "100110",
      "101011" when "100111",
      "000000" when "101000",
      "010110" when "101001",
      "001011" when "101010",
      "000000" when "101011",
      "101111" when "101100",
      "001100" when "101101",
      "101010" when "101110",
      "001110" when "101111",
      "000000" when "110000",
      "000000" when "110001",
      "100101" when "110010",
      "000000" when "110011",
      "011110" when "110100",
      "010001" when "110101",
      "000000" when "110110",
      "010111" when "110111",
      "001010" when "111000",
      "100001" when "111001",
      "100111" when "111010",
      "000000" when "111011",
      "100011" when "111100",
      "010011" when "111101",
      "000000" when "111110",
      "000101" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum1_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum1_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum1_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Sum1_2_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum1_2_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum12_2_impl_0_LUT_wIn_6_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum12_2_impl_0_LUT_wIn_6_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum12_2_impl_0_LUT_wIn_6_wOut_5 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "00000" when "000000",
      "00000" when "000001",
      "10001" when "000010",
      "00000" when "000011",
      "01111" when "000100",
      "00000" when "000101",
      "00000" when "000110",
      "00000" when "000111",
      "00000" when "001000",
      "01101" when "001001",
      "00000" when "001010",
      "00000" when "001011",
      "00100" when "001100",
      "00000" when "001101",
      "00000" when "001110",
      "00000" when "001111",
      "00000" when "010000",
      "00000" when "010001",
      "00000" when "010010",
      "00101" when "010011",
      "00011" when "010100",
      "00000" when "010101",
      "00000" when "010110",
      "00000" when "010111",
      "00000" when "011000",
      "00000" when "011001",
      "00000" when "011010",
      "00000" when "011011",
      "00000" when "011100",
      "00000" when "011101",
      "00000" when "011110",
      "00000" when "011111",
      "01001" when "100000",
      "00000" when "100001",
      "01010" when "100010",
      "00000" when "100011",
      "00000" when "100100",
      "00000" when "100101",
      "00000" when "100110",
      "10000" when "100111",
      "00000" when "101000",
      "00001" when "101001",
      "01000" when "101010",
      "00000" when "101011",
      "00000" when "101100",
      "00000" when "101101",
      "00000" when "101110",
      "00010" when "101111",
      "00000" when "110000",
      "00000" when "110001",
      "01011" when "110010",
      "00000" when "110011",
      "01100" when "110100",
      "10010" when "110101",
      "00000" when "110110",
      "00110" when "110111",
      "00000" when "111000",
      "00000" when "111001",
      "00000" when "111010",
      "00000" when "111011",
      "10011" when "111100",
      "00000" when "111101",
      "01110" when "111110",
      "00111" when "111111",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum12_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum12_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum12_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Sum12_2_impl_0_LUT_wIn_6_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum12_2_impl_0_LUT_wIn_6_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum12_2_impl_1_LUT_wIn_6_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum12_2_impl_1_LUT_wIn_6_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum12_2_impl_1_LUT_wIn_6_wOut_5 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "00000" when "000000",
      "00000" when "000001",
      "10010" when "000010",
      "00000" when "000011",
      "01100" when "000100",
      "00000" when "000101",
      "00000" when "000110",
      "00000" when "000111",
      "00000" when "001000",
      "01101" when "001001",
      "00000" when "001010",
      "00000" when "001011",
      "00011" when "001100",
      "00000" when "001101",
      "00000" when "001110",
      "00000" when "001111",
      "00000" when "010000",
      "00000" when "010001",
      "00000" when "010010",
      "00100" when "010011",
      "00010" when "010100",
      "00000" when "010101",
      "00000" when "010110",
      "00000" when "010111",
      "00000" when "011000",
      "01111" when "011001",
      "00000" when "011010",
      "00000" when "011011",
      "00000" when "011100",
      "00000" when "011101",
      "00000" when "011110",
      "00000" when "011111",
      "01000" when "100000",
      "00000" when "100001",
      "01001" when "100010",
      "00000" when "100011",
      "00000" when "100100",
      "00000" when "100101",
      "00000" when "100110",
      "01110" when "100111",
      "00000" when "101000",
      "00000" when "101001",
      "00111" when "101010",
      "00000" when "101011",
      "00000" when "101100",
      "00000" when "101101",
      "00000" when "101110",
      "00001" when "101111",
      "00000" when "110000",
      "00000" when "110001",
      "10011" when "110010",
      "00000" when "110011",
      "01010" when "110100",
      "10001" when "110101",
      "00000" when "110110",
      "00101" when "110111",
      "00000" when "111000",
      "00000" when "111001",
      "00000" when "111010",
      "00000" when "111011",
      "10000" when "111100",
      "00000" when "111101",
      "01011" when "111110",
      "00110" when "111111",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum12_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum12_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum12_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Sum12_2_impl_1_LUT_wIn_6_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum12_2_impl_1_LUT_wIn_6_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum15_2_impl_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum15_2_impl_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum15_2_impl_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "1010" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0100" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "1001" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0101" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0110" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0001" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "1011" when "100111",
      "0000" when "101000",
      "0010" when "101001",
      "0011" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "1000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0111" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "1100" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum15_2_impl_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum15_2_impl_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum15_2_impl_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Sum15_2_impl_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum15_2_impl_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum15_2_impl_1_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum15_2_impl_1_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum15_2_impl_1_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "1100" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0100" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "1011" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0101" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "1000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0001" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "1010" when "100111",
      "0000" when "101000",
      "0010" when "101001",
      "0011" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0111" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "1001" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0110" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum15_2_impl_1_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum15_2_impl_1_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum15_2_impl_1_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Sum15_2_impl_1_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum15_2_impl_1_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum2_2_impl_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum2_2_impl_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum2_2_impl_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "101" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "001" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "100" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "011" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "010" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum2_2_impl_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum2_2_impl_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum2_2_impl_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Sum2_2_impl_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum2_2_impl_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum2_2_impl_1_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum2_2_impl_1_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum2_2_impl_1_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "011" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "100" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "101" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "010" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "001" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum2_2_impl_1_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum2_2_impl_1_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum2_2_impl_1_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Sum2_2_impl_1_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum2_2_impl_1_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum26_1_impl_0_LUT_wIn_6_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum26_1_impl_0_LUT_wIn_6_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum26_1_impl_0_LUT_wIn_6_wOut_2 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "00" when "000000",
      "00" when "000001",
      "00" when "000010",
      "00" when "000011",
      "00" when "000100",
      "00" when "000101",
      "00" when "000110",
      "00" when "000111",
      "00" when "001000",
      "00" when "001001",
      "00" when "001010",
      "00" when "001011",
      "00" when "001100",
      "00" when "001101",
      "00" when "001110",
      "00" when "001111",
      "00" when "010000",
      "00" when "010001",
      "00" when "010010",
      "00" when "010011",
      "00" when "010100",
      "00" when "010101",
      "00" when "010110",
      "00" when "010111",
      "00" when "011000",
      "10" when "011001",
      "00" when "011010",
      "00" when "011011",
      "00" when "011100",
      "00" when "011101",
      "00" when "011110",
      "00" when "011111",
      "00" when "100000",
      "00" when "100001",
      "00" when "100010",
      "00" when "100011",
      "00" when "100100",
      "00" when "100101",
      "00" when "100110",
      "00" when "100111",
      "00" when "101000",
      "00" when "101001",
      "00" when "101010",
      "00" when "101011",
      "00" when "101100",
      "00" when "101101",
      "00" when "101110",
      "01" when "101111",
      "00" when "110000",
      "00" when "110001",
      "00" when "110010",
      "00" when "110011",
      "00" when "110100",
      "00" when "110101",
      "00" when "110110",
      "00" when "110111",
      "00" when "111000",
      "00" when "111001",
      "00" when "111010",
      "00" when "111011",
      "00" when "111100",
      "00" when "111101",
      "00" when "111110",
      "00" when "111111",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum26_1_impl_0_LUT_wIn_6_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum26_1_impl_0_LUT_wIn_6_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum26_1_impl_0_LUT_wIn_6_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Sum26_1_impl_0_LUT_wIn_6_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum26_1_impl_0_LUT_wIn_6_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum26_1_impl_1_LUT_wIn_6_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum26_1_impl_1_LUT_wIn_6_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum26_1_impl_1_LUT_wIn_6_wOut_2 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "00" when "000000",
      "00" when "000001",
      "00" when "000010",
      "00" when "000011",
      "00" when "000100",
      "00" when "000101",
      "00" when "000110",
      "00" when "000111",
      "00" when "001000",
      "00" when "001001",
      "00" when "001010",
      "00" when "001011",
      "00" when "001100",
      "00" when "001101",
      "00" when "001110",
      "00" when "001111",
      "00" when "010000",
      "00" when "010001",
      "00" when "010010",
      "00" when "010011",
      "00" when "010100",
      "00" when "010101",
      "00" when "010110",
      "00" when "010111",
      "00" when "011000",
      "10" when "011001",
      "00" when "011010",
      "00" when "011011",
      "00" when "011100",
      "00" when "011101",
      "00" when "011110",
      "00" when "011111",
      "00" when "100000",
      "00" when "100001",
      "00" when "100010",
      "00" when "100011",
      "00" when "100100",
      "00" when "100101",
      "00" when "100110",
      "00" when "100111",
      "00" when "101000",
      "00" when "101001",
      "00" when "101010",
      "00" when "101011",
      "00" when "101100",
      "00" when "101101",
      "00" when "101110",
      "01" when "101111",
      "00" when "110000",
      "00" when "110001",
      "00" when "110010",
      "00" when "110011",
      "00" when "110100",
      "00" when "110101",
      "00" when "110110",
      "00" when "110111",
      "00" when "111000",
      "00" when "111001",
      "00" when "111010",
      "00" when "111011",
      "00" when "111100",
      "00" when "111101",
      "00" when "111110",
      "00" when "111111",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum26_1_impl_1_LUT_wIn_6_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum26_1_impl_1_LUT_wIn_6_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum26_1_impl_1_LUT_wIn_6_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Sum26_1_impl_1_LUT_wIn_6_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum26_1_impl_1_LUT_wIn_6_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum41_2_impl_0_LUT_wIn_6_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum41_2_impl_0_LUT_wIn_6_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum41_2_impl_0_LUT_wIn_6_wOut_1 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0" when "000000",
      "0" when "000001",
      "0" when "000010",
      "0" when "000011",
      "0" when "000100",
      "0" when "000101",
      "0" when "000110",
      "0" when "000111",
      "0" when "001000",
      "0" when "001001",
      "0" when "001010",
      "0" when "001011",
      "0" when "001100",
      "0" when "001101",
      "0" when "001110",
      "0" when "001111",
      "0" when "010000",
      "0" when "010001",
      "0" when "010010",
      "0" when "010011",
      "0" when "010100",
      "0" when "010101",
      "0" when "010110",
      "0" when "010111",
      "0" when "011000",
      "0" when "011001",
      "0" when "011010",
      "0" when "011011",
      "0" when "011100",
      "0" when "011101",
      "0" when "011110",
      "0" when "011111",
      "0" when "100000",
      "0" when "100001",
      "0" when "100010",
      "0" when "100011",
      "0" when "100100",
      "0" when "100101",
      "0" when "100110",
      "0" when "100111",
      "0" when "101000",
      "0" when "101001",
      "0" when "101010",
      "0" when "101011",
      "0" when "101100",
      "0" when "101101",
      "0" when "101110",
      "1" when "101111",
      "0" when "110000",
      "0" when "110001",
      "0" when "110010",
      "0" when "110011",
      "0" when "110100",
      "0" when "110101",
      "0" when "110110",
      "0" when "110111",
      "0" when "111000",
      "0" when "111001",
      "0" when "111010",
      "0" when "111011",
      "0" when "111100",
      "0" when "111101",
      "0" when "111110",
      "0" when "111111",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum41_2_impl_0_LUT_wIn_6_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum41_2_impl_0_LUT_wIn_6_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum41_2_impl_0_LUT_wIn_6_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Sum41_2_impl_0_LUT_wIn_6_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum41_2_impl_0_LUT_wIn_6_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum41_2_impl_1_LUT_wIn_6_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum41_2_impl_1_LUT_wIn_6_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum41_2_impl_1_LUT_wIn_6_wOut_1 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0" when "000000",
      "0" when "000001",
      "0" when "000010",
      "0" when "000011",
      "0" when "000100",
      "0" when "000101",
      "0" when "000110",
      "0" when "000111",
      "0" when "001000",
      "0" when "001001",
      "0" when "001010",
      "0" when "001011",
      "0" when "001100",
      "0" when "001101",
      "0" when "001110",
      "0" when "001111",
      "0" when "010000",
      "0" when "010001",
      "0" when "010010",
      "0" when "010011",
      "0" when "010100",
      "0" when "010101",
      "0" when "010110",
      "0" when "010111",
      "0" when "011000",
      "0" when "011001",
      "0" when "011010",
      "0" when "011011",
      "0" when "011100",
      "0" when "011101",
      "0" when "011110",
      "0" when "011111",
      "0" when "100000",
      "0" when "100001",
      "0" when "100010",
      "0" when "100011",
      "0" when "100100",
      "0" when "100101",
      "0" when "100110",
      "0" when "100111",
      "0" when "101000",
      "0" when "101001",
      "0" when "101010",
      "0" when "101011",
      "0" when "101100",
      "0" when "101101",
      "0" when "101110",
      "1" when "101111",
      "0" when "110000",
      "0" when "110001",
      "0" when "110010",
      "0" when "110011",
      "0" when "110100",
      "0" when "110101",
      "0" when "110110",
      "0" when "110111",
      "0" when "111000",
      "0" when "111001",
      "0" when "111010",
      "0" when "111011",
      "0" when "111100",
      "0" when "111101",
      "0" when "111110",
      "0" when "111111",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum41_2_impl_1_LUT_wIn_6_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum41_2_impl_1_LUT_wIn_6_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum41_2_impl_1_LUT_wIn_6_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Sum41_2_impl_1_LUT_wIn_6_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum41_2_impl_1_LUT_wIn_6_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum42_2_impl_0_LUT_wIn_6_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum42_2_impl_0_LUT_wIn_6_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum42_2_impl_0_LUT_wIn_6_wOut_1 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0" when "000000",
      "0" when "000001",
      "0" when "000010",
      "0" when "000011",
      "0" when "000100",
      "0" when "000101",
      "0" when "000110",
      "0" when "000111",
      "0" when "001000",
      "0" when "001001",
      "0" when "001010",
      "0" when "001011",
      "0" when "001100",
      "0" when "001101",
      "0" when "001110",
      "0" when "001111",
      "0" when "010000",
      "0" when "010001",
      "0" when "010010",
      "0" when "010011",
      "0" when "010100",
      "0" when "010101",
      "0" when "010110",
      "0" when "010111",
      "0" when "011000",
      "0" when "011001",
      "0" when "011010",
      "0" when "011011",
      "0" when "011100",
      "0" when "011101",
      "0" when "011110",
      "0" when "011111",
      "0" when "100000",
      "0" when "100001",
      "0" when "100010",
      "0" when "100011",
      "0" when "100100",
      "0" when "100101",
      "0" when "100110",
      "0" when "100111",
      "0" when "101000",
      "0" when "101001",
      "0" when "101010",
      "0" when "101011",
      "0" when "101100",
      "0" when "101101",
      "0" when "101110",
      "1" when "101111",
      "0" when "110000",
      "0" when "110001",
      "0" when "110010",
      "0" when "110011",
      "0" when "110100",
      "0" when "110101",
      "0" when "110110",
      "0" when "110111",
      "0" when "111000",
      "0" when "111001",
      "0" when "111010",
      "0" when "111011",
      "0" when "111100",
      "0" when "111101",
      "0" when "111110",
      "0" when "111111",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum42_2_impl_0_LUT_wIn_6_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum42_2_impl_0_LUT_wIn_6_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum42_2_impl_0_LUT_wIn_6_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Sum42_2_impl_0_LUT_wIn_6_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum42_2_impl_0_LUT_wIn_6_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Sum42_2_impl_1_LUT_wIn_6_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum42_2_impl_1_LUT_wIn_6_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum42_2_impl_1_LUT_wIn_6_wOut_1 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0" when "000000",
      "0" when "000001",
      "0" when "000010",
      "0" when "000011",
      "1" when "000100",
      "0" when "000101",
      "0" when "000110",
      "0" when "000111",
      "0" when "001000",
      "0" when "001001",
      "0" when "001010",
      "0" when "001011",
      "0" when "001100",
      "0" when "001101",
      "0" when "001110",
      "0" when "001111",
      "0" when "010000",
      "0" when "010001",
      "0" when "010010",
      "0" when "010011",
      "0" when "010100",
      "0" when "010101",
      "0" when "010110",
      "0" when "010111",
      "0" when "011000",
      "0" when "011001",
      "0" when "011010",
      "0" when "011011",
      "0" when "011100",
      "0" when "011101",
      "0" when "011110",
      "0" when "011111",
      "0" when "100000",
      "0" when "100001",
      "0" when "100010",
      "0" when "100011",
      "0" when "100100",
      "0" when "100101",
      "0" when "100110",
      "0" when "100111",
      "0" when "101000",
      "0" when "101001",
      "0" when "101010",
      "0" when "101011",
      "0" when "101100",
      "0" when "101101",
      "0" when "101110",
      "0" when "101111",
      "0" when "110000",
      "0" when "110001",
      "0" when "110010",
      "0" when "110011",
      "0" when "110100",
      "0" when "110101",
      "0" when "110110",
      "0" when "110111",
      "0" when "111000",
      "0" when "111001",
      "0" when "111010",
      "0" when "111011",
      "0" when "111100",
      "0" when "111101",
      "0" when "111110",
      "0" when "111111",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Sum42_2_impl_1_LUT_wIn_6_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Sum42_2_impl_1_LUT_wIn_6_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Sum42_2_impl_1_LUT_wIn_6_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Sum42_2_impl_1_LUT_wIn_6_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Sum42_2_impl_1_LUT_wIn_6_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--              GenericLut_LUTData_MUX_Out2_0_0_LUT_wIn_6_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Out2_0_0_LUT_wIn_6_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Out2_0_0_LUT_wIn_6_wOut_2 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "00" when "000000",
      "01" when "000001",
      "00" when "000010",
      "00" when "000011",
      "00" when "000100",
      "00" when "000101",
      "00" when "000110",
      "00" when "000111",
      "00" when "001000",
      "00" when "001001",
      "00" when "001010",
      "00" when "001011",
      "00" when "001100",
      "00" when "001101",
      "00" when "001110",
      "00" when "001111",
      "00" when "010000",
      "00" when "010001",
      "00" when "010010",
      "00" when "010011",
      "00" when "010100",
      "00" when "010101",
      "00" when "010110",
      "10" when "010111",
      "00" when "011000",
      "00" when "011001",
      "00" when "011010",
      "00" when "011011",
      "00" when "011100",
      "00" when "011101",
      "00" when "011110",
      "00" when "011111",
      "00" when "100000",
      "00" when "100001",
      "00" when "100010",
      "00" when "100011",
      "00" when "100100",
      "00" when "100101",
      "00" when "100110",
      "00" when "100111",
      "00" when "101000",
      "00" when "101001",
      "00" when "101010",
      "00" when "101011",
      "00" when "101100",
      "00" when "101101",
      "00" when "101110",
      "00" when "101111",
      "00" when "110000",
      "00" when "110001",
      "00" when "110010",
      "00" when "110011",
      "00" when "110100",
      "00" when "110101",
      "00" when "110110",
      "00" when "110111",
      "00" when "111000",
      "00" when "111001",
      "00" when "111010",
      "00" when "111011",
      "00" when "111100",
      "00" when "111101",
      "00" when "111110",
      "00" when "111111",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--     GenericLut_LUTData_MUX_Out2_0_0_LUT_wIn_6_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Out2_0_0_LUT_wIn_6_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Out2_0_0_LUT_wIn_6_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Out2_0_0_LUT_wIn_6_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Out2_0_0_LUT_wIn_6_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 68 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      Y <= s67;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      Y <= s15;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      Y <= s18;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 24 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      Y <= s23;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 53 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      Y <= s52;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_100_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 100 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_100_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_100_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      Y <= s99;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_684_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 684 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_684_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_684_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
signal s558 : std_logic_vector(33 downto 0) := (others => '0');
signal s559 : std_logic_vector(33 downto 0) := (others => '0');
signal s560 : std_logic_vector(33 downto 0) := (others => '0');
signal s561 : std_logic_vector(33 downto 0) := (others => '0');
signal s562 : std_logic_vector(33 downto 0) := (others => '0');
signal s563 : std_logic_vector(33 downto 0) := (others => '0');
signal s564 : std_logic_vector(33 downto 0) := (others => '0');
signal s565 : std_logic_vector(33 downto 0) := (others => '0');
signal s566 : std_logic_vector(33 downto 0) := (others => '0');
signal s567 : std_logic_vector(33 downto 0) := (others => '0');
signal s568 : std_logic_vector(33 downto 0) := (others => '0');
signal s569 : std_logic_vector(33 downto 0) := (others => '0');
signal s570 : std_logic_vector(33 downto 0) := (others => '0');
signal s571 : std_logic_vector(33 downto 0) := (others => '0');
signal s572 : std_logic_vector(33 downto 0) := (others => '0');
signal s573 : std_logic_vector(33 downto 0) := (others => '0');
signal s574 : std_logic_vector(33 downto 0) := (others => '0');
signal s575 : std_logic_vector(33 downto 0) := (others => '0');
signal s576 : std_logic_vector(33 downto 0) := (others => '0');
signal s577 : std_logic_vector(33 downto 0) := (others => '0');
signal s578 : std_logic_vector(33 downto 0) := (others => '0');
signal s579 : std_logic_vector(33 downto 0) := (others => '0');
signal s580 : std_logic_vector(33 downto 0) := (others => '0');
signal s581 : std_logic_vector(33 downto 0) := (others => '0');
signal s582 : std_logic_vector(33 downto 0) := (others => '0');
signal s583 : std_logic_vector(33 downto 0) := (others => '0');
signal s584 : std_logic_vector(33 downto 0) := (others => '0');
signal s585 : std_logic_vector(33 downto 0) := (others => '0');
signal s586 : std_logic_vector(33 downto 0) := (others => '0');
signal s587 : std_logic_vector(33 downto 0) := (others => '0');
signal s588 : std_logic_vector(33 downto 0) := (others => '0');
signal s589 : std_logic_vector(33 downto 0) := (others => '0');
signal s590 : std_logic_vector(33 downto 0) := (others => '0');
signal s591 : std_logic_vector(33 downto 0) := (others => '0');
signal s592 : std_logic_vector(33 downto 0) := (others => '0');
signal s593 : std_logic_vector(33 downto 0) := (others => '0');
signal s594 : std_logic_vector(33 downto 0) := (others => '0');
signal s595 : std_logic_vector(33 downto 0) := (others => '0');
signal s596 : std_logic_vector(33 downto 0) := (others => '0');
signal s597 : std_logic_vector(33 downto 0) := (others => '0');
signal s598 : std_logic_vector(33 downto 0) := (others => '0');
signal s599 : std_logic_vector(33 downto 0) := (others => '0');
signal s600 : std_logic_vector(33 downto 0) := (others => '0');
signal s601 : std_logic_vector(33 downto 0) := (others => '0');
signal s602 : std_logic_vector(33 downto 0) := (others => '0');
signal s603 : std_logic_vector(33 downto 0) := (others => '0');
signal s604 : std_logic_vector(33 downto 0) := (others => '0');
signal s605 : std_logic_vector(33 downto 0) := (others => '0');
signal s606 : std_logic_vector(33 downto 0) := (others => '0');
signal s607 : std_logic_vector(33 downto 0) := (others => '0');
signal s608 : std_logic_vector(33 downto 0) := (others => '0');
signal s609 : std_logic_vector(33 downto 0) := (others => '0');
signal s610 : std_logic_vector(33 downto 0) := (others => '0');
signal s611 : std_logic_vector(33 downto 0) := (others => '0');
signal s612 : std_logic_vector(33 downto 0) := (others => '0');
signal s613 : std_logic_vector(33 downto 0) := (others => '0');
signal s614 : std_logic_vector(33 downto 0) := (others => '0');
signal s615 : std_logic_vector(33 downto 0) := (others => '0');
signal s616 : std_logic_vector(33 downto 0) := (others => '0');
signal s617 : std_logic_vector(33 downto 0) := (others => '0');
signal s618 : std_logic_vector(33 downto 0) := (others => '0');
signal s619 : std_logic_vector(33 downto 0) := (others => '0');
signal s620 : std_logic_vector(33 downto 0) := (others => '0');
signal s621 : std_logic_vector(33 downto 0) := (others => '0');
signal s622 : std_logic_vector(33 downto 0) := (others => '0');
signal s623 : std_logic_vector(33 downto 0) := (others => '0');
signal s624 : std_logic_vector(33 downto 0) := (others => '0');
signal s625 : std_logic_vector(33 downto 0) := (others => '0');
signal s626 : std_logic_vector(33 downto 0) := (others => '0');
signal s627 : std_logic_vector(33 downto 0) := (others => '0');
signal s628 : std_logic_vector(33 downto 0) := (others => '0');
signal s629 : std_logic_vector(33 downto 0) := (others => '0');
signal s630 : std_logic_vector(33 downto 0) := (others => '0');
signal s631 : std_logic_vector(33 downto 0) := (others => '0');
signal s632 : std_logic_vector(33 downto 0) := (others => '0');
signal s633 : std_logic_vector(33 downto 0) := (others => '0');
signal s634 : std_logic_vector(33 downto 0) := (others => '0');
signal s635 : std_logic_vector(33 downto 0) := (others => '0');
signal s636 : std_logic_vector(33 downto 0) := (others => '0');
signal s637 : std_logic_vector(33 downto 0) := (others => '0');
signal s638 : std_logic_vector(33 downto 0) := (others => '0');
signal s639 : std_logic_vector(33 downto 0) := (others => '0');
signal s640 : std_logic_vector(33 downto 0) := (others => '0');
signal s641 : std_logic_vector(33 downto 0) := (others => '0');
signal s642 : std_logic_vector(33 downto 0) := (others => '0');
signal s643 : std_logic_vector(33 downto 0) := (others => '0');
signal s644 : std_logic_vector(33 downto 0) := (others => '0');
signal s645 : std_logic_vector(33 downto 0) := (others => '0');
signal s646 : std_logic_vector(33 downto 0) := (others => '0');
signal s647 : std_logic_vector(33 downto 0) := (others => '0');
signal s648 : std_logic_vector(33 downto 0) := (others => '0');
signal s649 : std_logic_vector(33 downto 0) := (others => '0');
signal s650 : std_logic_vector(33 downto 0) := (others => '0');
signal s651 : std_logic_vector(33 downto 0) := (others => '0');
signal s652 : std_logic_vector(33 downto 0) := (others => '0');
signal s653 : std_logic_vector(33 downto 0) := (others => '0');
signal s654 : std_logic_vector(33 downto 0) := (others => '0');
signal s655 : std_logic_vector(33 downto 0) := (others => '0');
signal s656 : std_logic_vector(33 downto 0) := (others => '0');
signal s657 : std_logic_vector(33 downto 0) := (others => '0');
signal s658 : std_logic_vector(33 downto 0) := (others => '0');
signal s659 : std_logic_vector(33 downto 0) := (others => '0');
signal s660 : std_logic_vector(33 downto 0) := (others => '0');
signal s661 : std_logic_vector(33 downto 0) := (others => '0');
signal s662 : std_logic_vector(33 downto 0) := (others => '0');
signal s663 : std_logic_vector(33 downto 0) := (others => '0');
signal s664 : std_logic_vector(33 downto 0) := (others => '0');
signal s665 : std_logic_vector(33 downto 0) := (others => '0');
signal s666 : std_logic_vector(33 downto 0) := (others => '0');
signal s667 : std_logic_vector(33 downto 0) := (others => '0');
signal s668 : std_logic_vector(33 downto 0) := (others => '0');
signal s669 : std_logic_vector(33 downto 0) := (others => '0');
signal s670 : std_logic_vector(33 downto 0) := (others => '0');
signal s671 : std_logic_vector(33 downto 0) := (others => '0');
signal s672 : std_logic_vector(33 downto 0) := (others => '0');
signal s673 : std_logic_vector(33 downto 0) := (others => '0');
signal s674 : std_logic_vector(33 downto 0) := (others => '0');
signal s675 : std_logic_vector(33 downto 0) := (others => '0');
signal s676 : std_logic_vector(33 downto 0) := (others => '0');
signal s677 : std_logic_vector(33 downto 0) := (others => '0');
signal s678 : std_logic_vector(33 downto 0) := (others => '0');
signal s679 : std_logic_vector(33 downto 0) := (others => '0');
signal s680 : std_logic_vector(33 downto 0) := (others => '0');
signal s681 : std_logic_vector(33 downto 0) := (others => '0');
signal s682 : std_logic_vector(33 downto 0) := (others => '0');
signal s683 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
      s558 <= "0000000000000000000000000000000000";
      s559 <= "0000000000000000000000000000000000";
      s560 <= "0000000000000000000000000000000000";
      s561 <= "0000000000000000000000000000000000";
      s562 <= "0000000000000000000000000000000000";
      s563 <= "0000000000000000000000000000000000";
      s564 <= "0000000000000000000000000000000000";
      s565 <= "0000000000000000000000000000000000";
      s566 <= "0000000000000000000000000000000000";
      s567 <= "0000000000000000000000000000000000";
      s568 <= "0000000000000000000000000000000000";
      s569 <= "0000000000000000000000000000000000";
      s570 <= "0000000000000000000000000000000000";
      s571 <= "0000000000000000000000000000000000";
      s572 <= "0000000000000000000000000000000000";
      s573 <= "0000000000000000000000000000000000";
      s574 <= "0000000000000000000000000000000000";
      s575 <= "0000000000000000000000000000000000";
      s576 <= "0000000000000000000000000000000000";
      s577 <= "0000000000000000000000000000000000";
      s578 <= "0000000000000000000000000000000000";
      s579 <= "0000000000000000000000000000000000";
      s580 <= "0000000000000000000000000000000000";
      s581 <= "0000000000000000000000000000000000";
      s582 <= "0000000000000000000000000000000000";
      s583 <= "0000000000000000000000000000000000";
      s584 <= "0000000000000000000000000000000000";
      s585 <= "0000000000000000000000000000000000";
      s586 <= "0000000000000000000000000000000000";
      s587 <= "0000000000000000000000000000000000";
      s588 <= "0000000000000000000000000000000000";
      s589 <= "0000000000000000000000000000000000";
      s590 <= "0000000000000000000000000000000000";
      s591 <= "0000000000000000000000000000000000";
      s592 <= "0000000000000000000000000000000000";
      s593 <= "0000000000000000000000000000000000";
      s594 <= "0000000000000000000000000000000000";
      s595 <= "0000000000000000000000000000000000";
      s596 <= "0000000000000000000000000000000000";
      s597 <= "0000000000000000000000000000000000";
      s598 <= "0000000000000000000000000000000000";
      s599 <= "0000000000000000000000000000000000";
      s600 <= "0000000000000000000000000000000000";
      s601 <= "0000000000000000000000000000000000";
      s602 <= "0000000000000000000000000000000000";
      s603 <= "0000000000000000000000000000000000";
      s604 <= "0000000000000000000000000000000000";
      s605 <= "0000000000000000000000000000000000";
      s606 <= "0000000000000000000000000000000000";
      s607 <= "0000000000000000000000000000000000";
      s608 <= "0000000000000000000000000000000000";
      s609 <= "0000000000000000000000000000000000";
      s610 <= "0000000000000000000000000000000000";
      s611 <= "0000000000000000000000000000000000";
      s612 <= "0000000000000000000000000000000000";
      s613 <= "0000000000000000000000000000000000";
      s614 <= "0000000000000000000000000000000000";
      s615 <= "0000000000000000000000000000000000";
      s616 <= "0000000000000000000000000000000000";
      s617 <= "0000000000000000000000000000000000";
      s618 <= "0000000000000000000000000000000000";
      s619 <= "0000000000000000000000000000000000";
      s620 <= "0000000000000000000000000000000000";
      s621 <= "0000000000000000000000000000000000";
      s622 <= "0000000000000000000000000000000000";
      s623 <= "0000000000000000000000000000000000";
      s624 <= "0000000000000000000000000000000000";
      s625 <= "0000000000000000000000000000000000";
      s626 <= "0000000000000000000000000000000000";
      s627 <= "0000000000000000000000000000000000";
      s628 <= "0000000000000000000000000000000000";
      s629 <= "0000000000000000000000000000000000";
      s630 <= "0000000000000000000000000000000000";
      s631 <= "0000000000000000000000000000000000";
      s632 <= "0000000000000000000000000000000000";
      s633 <= "0000000000000000000000000000000000";
      s634 <= "0000000000000000000000000000000000";
      s635 <= "0000000000000000000000000000000000";
      s636 <= "0000000000000000000000000000000000";
      s637 <= "0000000000000000000000000000000000";
      s638 <= "0000000000000000000000000000000000";
      s639 <= "0000000000000000000000000000000000";
      s640 <= "0000000000000000000000000000000000";
      s641 <= "0000000000000000000000000000000000";
      s642 <= "0000000000000000000000000000000000";
      s643 <= "0000000000000000000000000000000000";
      s644 <= "0000000000000000000000000000000000";
      s645 <= "0000000000000000000000000000000000";
      s646 <= "0000000000000000000000000000000000";
      s647 <= "0000000000000000000000000000000000";
      s648 <= "0000000000000000000000000000000000";
      s649 <= "0000000000000000000000000000000000";
      s650 <= "0000000000000000000000000000000000";
      s651 <= "0000000000000000000000000000000000";
      s652 <= "0000000000000000000000000000000000";
      s653 <= "0000000000000000000000000000000000";
      s654 <= "0000000000000000000000000000000000";
      s655 <= "0000000000000000000000000000000000";
      s656 <= "0000000000000000000000000000000000";
      s657 <= "0000000000000000000000000000000000";
      s658 <= "0000000000000000000000000000000000";
      s659 <= "0000000000000000000000000000000000";
      s660 <= "0000000000000000000000000000000000";
      s661 <= "0000000000000000000000000000000000";
      s662 <= "0000000000000000000000000000000000";
      s663 <= "0000000000000000000000000000000000";
      s664 <= "0000000000000000000000000000000000";
      s665 <= "0000000000000000000000000000000000";
      s666 <= "0000000000000000000000000000000000";
      s667 <= "0000000000000000000000000000000000";
      s668 <= "0000000000000000000000000000000000";
      s669 <= "0000000000000000000000000000000000";
      s670 <= "0000000000000000000000000000000000";
      s671 <= "0000000000000000000000000000000000";
      s672 <= "0000000000000000000000000000000000";
      s673 <= "0000000000000000000000000000000000";
      s674 <= "0000000000000000000000000000000000";
      s675 <= "0000000000000000000000000000000000";
      s676 <= "0000000000000000000000000000000000";
      s677 <= "0000000000000000000000000000000000";
      s678 <= "0000000000000000000000000000000000";
      s679 <= "0000000000000000000000000000000000";
      s680 <= "0000000000000000000000000000000000";
      s681 <= "0000000000000000000000000000000000";
      s682 <= "0000000000000000000000000000000000";
      s683 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      s558 <= s557;
      s559 <= s558;
      s560 <= s559;
      s561 <= s560;
      s562 <= s561;
      s563 <= s562;
      s564 <= s563;
      s565 <= s564;
      s566 <= s565;
      s567 <= s566;
      s568 <= s567;
      s569 <= s568;
      s570 <= s569;
      s571 <= s570;
      s572 <= s571;
      s573 <= s572;
      s574 <= s573;
      s575 <= s574;
      s576 <= s575;
      s577 <= s576;
      s578 <= s577;
      s579 <= s578;
      s580 <= s579;
      s581 <= s580;
      s582 <= s581;
      s583 <= s582;
      s584 <= s583;
      s585 <= s584;
      s586 <= s585;
      s587 <= s586;
      s588 <= s587;
      s589 <= s588;
      s590 <= s589;
      s591 <= s590;
      s592 <= s591;
      s593 <= s592;
      s594 <= s593;
      s595 <= s594;
      s596 <= s595;
      s597 <= s596;
      s598 <= s597;
      s599 <= s598;
      s600 <= s599;
      s601 <= s600;
      s602 <= s601;
      s603 <= s602;
      s604 <= s603;
      s605 <= s604;
      s606 <= s605;
      s607 <= s606;
      s608 <= s607;
      s609 <= s608;
      s610 <= s609;
      s611 <= s610;
      s612 <= s611;
      s613 <= s612;
      s614 <= s613;
      s615 <= s614;
      s616 <= s615;
      s617 <= s616;
      s618 <= s617;
      s619 <= s618;
      s620 <= s619;
      s621 <= s620;
      s622 <= s621;
      s623 <= s622;
      s624 <= s623;
      s625 <= s624;
      s626 <= s625;
      s627 <= s626;
      s628 <= s627;
      s629 <= s628;
      s630 <= s629;
      s631 <= s630;
      s632 <= s631;
      s633 <= s632;
      s634 <= s633;
      s635 <= s634;
      s636 <= s635;
      s637 <= s636;
      s638 <= s637;
      s639 <= s638;
      s640 <= s639;
      s641 <= s640;
      s642 <= s641;
      s643 <= s642;
      s644 <= s643;
      s645 <= s644;
      s646 <= s645;
      s647 <= s646;
      s648 <= s647;
      s649 <= s648;
      s650 <= s649;
      s651 <= s650;
      s652 <= s651;
      s653 <= s652;
      s654 <= s653;
      s655 <= s654;
      s656 <= s655;
      s657 <= s656;
      s658 <= s657;
      s659 <= s658;
      s660 <= s659;
      s661 <= s660;
      s662 <= s661;
      s663 <= s662;
      s664 <= s663;
      s665 <= s664;
      s666 <= s665;
      s667 <= s666;
      s668 <= s667;
      s669 <= s668;
      s670 <= s669;
      s671 <= s670;
      s672 <= s671;
      s673 <= s672;
      s674 <= s673;
      s675 <= s674;
      s676 <= s675;
      s677 <= s676;
      s678 <= s677;
      s679 <= s678;
      s680 <= s679;
      s681 <= s680;
      s682 <= s681;
      s683 <= s682;
      Y <= s683;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_746_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 746 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_746_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_746_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
signal s558 : std_logic_vector(33 downto 0) := (others => '0');
signal s559 : std_logic_vector(33 downto 0) := (others => '0');
signal s560 : std_logic_vector(33 downto 0) := (others => '0');
signal s561 : std_logic_vector(33 downto 0) := (others => '0');
signal s562 : std_logic_vector(33 downto 0) := (others => '0');
signal s563 : std_logic_vector(33 downto 0) := (others => '0');
signal s564 : std_logic_vector(33 downto 0) := (others => '0');
signal s565 : std_logic_vector(33 downto 0) := (others => '0');
signal s566 : std_logic_vector(33 downto 0) := (others => '0');
signal s567 : std_logic_vector(33 downto 0) := (others => '0');
signal s568 : std_logic_vector(33 downto 0) := (others => '0');
signal s569 : std_logic_vector(33 downto 0) := (others => '0');
signal s570 : std_logic_vector(33 downto 0) := (others => '0');
signal s571 : std_logic_vector(33 downto 0) := (others => '0');
signal s572 : std_logic_vector(33 downto 0) := (others => '0');
signal s573 : std_logic_vector(33 downto 0) := (others => '0');
signal s574 : std_logic_vector(33 downto 0) := (others => '0');
signal s575 : std_logic_vector(33 downto 0) := (others => '0');
signal s576 : std_logic_vector(33 downto 0) := (others => '0');
signal s577 : std_logic_vector(33 downto 0) := (others => '0');
signal s578 : std_logic_vector(33 downto 0) := (others => '0');
signal s579 : std_logic_vector(33 downto 0) := (others => '0');
signal s580 : std_logic_vector(33 downto 0) := (others => '0');
signal s581 : std_logic_vector(33 downto 0) := (others => '0');
signal s582 : std_logic_vector(33 downto 0) := (others => '0');
signal s583 : std_logic_vector(33 downto 0) := (others => '0');
signal s584 : std_logic_vector(33 downto 0) := (others => '0');
signal s585 : std_logic_vector(33 downto 0) := (others => '0');
signal s586 : std_logic_vector(33 downto 0) := (others => '0');
signal s587 : std_logic_vector(33 downto 0) := (others => '0');
signal s588 : std_logic_vector(33 downto 0) := (others => '0');
signal s589 : std_logic_vector(33 downto 0) := (others => '0');
signal s590 : std_logic_vector(33 downto 0) := (others => '0');
signal s591 : std_logic_vector(33 downto 0) := (others => '0');
signal s592 : std_logic_vector(33 downto 0) := (others => '0');
signal s593 : std_logic_vector(33 downto 0) := (others => '0');
signal s594 : std_logic_vector(33 downto 0) := (others => '0');
signal s595 : std_logic_vector(33 downto 0) := (others => '0');
signal s596 : std_logic_vector(33 downto 0) := (others => '0');
signal s597 : std_logic_vector(33 downto 0) := (others => '0');
signal s598 : std_logic_vector(33 downto 0) := (others => '0');
signal s599 : std_logic_vector(33 downto 0) := (others => '0');
signal s600 : std_logic_vector(33 downto 0) := (others => '0');
signal s601 : std_logic_vector(33 downto 0) := (others => '0');
signal s602 : std_logic_vector(33 downto 0) := (others => '0');
signal s603 : std_logic_vector(33 downto 0) := (others => '0');
signal s604 : std_logic_vector(33 downto 0) := (others => '0');
signal s605 : std_logic_vector(33 downto 0) := (others => '0');
signal s606 : std_logic_vector(33 downto 0) := (others => '0');
signal s607 : std_logic_vector(33 downto 0) := (others => '0');
signal s608 : std_logic_vector(33 downto 0) := (others => '0');
signal s609 : std_logic_vector(33 downto 0) := (others => '0');
signal s610 : std_logic_vector(33 downto 0) := (others => '0');
signal s611 : std_logic_vector(33 downto 0) := (others => '0');
signal s612 : std_logic_vector(33 downto 0) := (others => '0');
signal s613 : std_logic_vector(33 downto 0) := (others => '0');
signal s614 : std_logic_vector(33 downto 0) := (others => '0');
signal s615 : std_logic_vector(33 downto 0) := (others => '0');
signal s616 : std_logic_vector(33 downto 0) := (others => '0');
signal s617 : std_logic_vector(33 downto 0) := (others => '0');
signal s618 : std_logic_vector(33 downto 0) := (others => '0');
signal s619 : std_logic_vector(33 downto 0) := (others => '0');
signal s620 : std_logic_vector(33 downto 0) := (others => '0');
signal s621 : std_logic_vector(33 downto 0) := (others => '0');
signal s622 : std_logic_vector(33 downto 0) := (others => '0');
signal s623 : std_logic_vector(33 downto 0) := (others => '0');
signal s624 : std_logic_vector(33 downto 0) := (others => '0');
signal s625 : std_logic_vector(33 downto 0) := (others => '0');
signal s626 : std_logic_vector(33 downto 0) := (others => '0');
signal s627 : std_logic_vector(33 downto 0) := (others => '0');
signal s628 : std_logic_vector(33 downto 0) := (others => '0');
signal s629 : std_logic_vector(33 downto 0) := (others => '0');
signal s630 : std_logic_vector(33 downto 0) := (others => '0');
signal s631 : std_logic_vector(33 downto 0) := (others => '0');
signal s632 : std_logic_vector(33 downto 0) := (others => '0');
signal s633 : std_logic_vector(33 downto 0) := (others => '0');
signal s634 : std_logic_vector(33 downto 0) := (others => '0');
signal s635 : std_logic_vector(33 downto 0) := (others => '0');
signal s636 : std_logic_vector(33 downto 0) := (others => '0');
signal s637 : std_logic_vector(33 downto 0) := (others => '0');
signal s638 : std_logic_vector(33 downto 0) := (others => '0');
signal s639 : std_logic_vector(33 downto 0) := (others => '0');
signal s640 : std_logic_vector(33 downto 0) := (others => '0');
signal s641 : std_logic_vector(33 downto 0) := (others => '0');
signal s642 : std_logic_vector(33 downto 0) := (others => '0');
signal s643 : std_logic_vector(33 downto 0) := (others => '0');
signal s644 : std_logic_vector(33 downto 0) := (others => '0');
signal s645 : std_logic_vector(33 downto 0) := (others => '0');
signal s646 : std_logic_vector(33 downto 0) := (others => '0');
signal s647 : std_logic_vector(33 downto 0) := (others => '0');
signal s648 : std_logic_vector(33 downto 0) := (others => '0');
signal s649 : std_logic_vector(33 downto 0) := (others => '0');
signal s650 : std_logic_vector(33 downto 0) := (others => '0');
signal s651 : std_logic_vector(33 downto 0) := (others => '0');
signal s652 : std_logic_vector(33 downto 0) := (others => '0');
signal s653 : std_logic_vector(33 downto 0) := (others => '0');
signal s654 : std_logic_vector(33 downto 0) := (others => '0');
signal s655 : std_logic_vector(33 downto 0) := (others => '0');
signal s656 : std_logic_vector(33 downto 0) := (others => '0');
signal s657 : std_logic_vector(33 downto 0) := (others => '0');
signal s658 : std_logic_vector(33 downto 0) := (others => '0');
signal s659 : std_logic_vector(33 downto 0) := (others => '0');
signal s660 : std_logic_vector(33 downto 0) := (others => '0');
signal s661 : std_logic_vector(33 downto 0) := (others => '0');
signal s662 : std_logic_vector(33 downto 0) := (others => '0');
signal s663 : std_logic_vector(33 downto 0) := (others => '0');
signal s664 : std_logic_vector(33 downto 0) := (others => '0');
signal s665 : std_logic_vector(33 downto 0) := (others => '0');
signal s666 : std_logic_vector(33 downto 0) := (others => '0');
signal s667 : std_logic_vector(33 downto 0) := (others => '0');
signal s668 : std_logic_vector(33 downto 0) := (others => '0');
signal s669 : std_logic_vector(33 downto 0) := (others => '0');
signal s670 : std_logic_vector(33 downto 0) := (others => '0');
signal s671 : std_logic_vector(33 downto 0) := (others => '0');
signal s672 : std_logic_vector(33 downto 0) := (others => '0');
signal s673 : std_logic_vector(33 downto 0) := (others => '0');
signal s674 : std_logic_vector(33 downto 0) := (others => '0');
signal s675 : std_logic_vector(33 downto 0) := (others => '0');
signal s676 : std_logic_vector(33 downto 0) := (others => '0');
signal s677 : std_logic_vector(33 downto 0) := (others => '0');
signal s678 : std_logic_vector(33 downto 0) := (others => '0');
signal s679 : std_logic_vector(33 downto 0) := (others => '0');
signal s680 : std_logic_vector(33 downto 0) := (others => '0');
signal s681 : std_logic_vector(33 downto 0) := (others => '0');
signal s682 : std_logic_vector(33 downto 0) := (others => '0');
signal s683 : std_logic_vector(33 downto 0) := (others => '0');
signal s684 : std_logic_vector(33 downto 0) := (others => '0');
signal s685 : std_logic_vector(33 downto 0) := (others => '0');
signal s686 : std_logic_vector(33 downto 0) := (others => '0');
signal s687 : std_logic_vector(33 downto 0) := (others => '0');
signal s688 : std_logic_vector(33 downto 0) := (others => '0');
signal s689 : std_logic_vector(33 downto 0) := (others => '0');
signal s690 : std_logic_vector(33 downto 0) := (others => '0');
signal s691 : std_logic_vector(33 downto 0) := (others => '0');
signal s692 : std_logic_vector(33 downto 0) := (others => '0');
signal s693 : std_logic_vector(33 downto 0) := (others => '0');
signal s694 : std_logic_vector(33 downto 0) := (others => '0');
signal s695 : std_logic_vector(33 downto 0) := (others => '0');
signal s696 : std_logic_vector(33 downto 0) := (others => '0');
signal s697 : std_logic_vector(33 downto 0) := (others => '0');
signal s698 : std_logic_vector(33 downto 0) := (others => '0');
signal s699 : std_logic_vector(33 downto 0) := (others => '0');
signal s700 : std_logic_vector(33 downto 0) := (others => '0');
signal s701 : std_logic_vector(33 downto 0) := (others => '0');
signal s702 : std_logic_vector(33 downto 0) := (others => '0');
signal s703 : std_logic_vector(33 downto 0) := (others => '0');
signal s704 : std_logic_vector(33 downto 0) := (others => '0');
signal s705 : std_logic_vector(33 downto 0) := (others => '0');
signal s706 : std_logic_vector(33 downto 0) := (others => '0');
signal s707 : std_logic_vector(33 downto 0) := (others => '0');
signal s708 : std_logic_vector(33 downto 0) := (others => '0');
signal s709 : std_logic_vector(33 downto 0) := (others => '0');
signal s710 : std_logic_vector(33 downto 0) := (others => '0');
signal s711 : std_logic_vector(33 downto 0) := (others => '0');
signal s712 : std_logic_vector(33 downto 0) := (others => '0');
signal s713 : std_logic_vector(33 downto 0) := (others => '0');
signal s714 : std_logic_vector(33 downto 0) := (others => '0');
signal s715 : std_logic_vector(33 downto 0) := (others => '0');
signal s716 : std_logic_vector(33 downto 0) := (others => '0');
signal s717 : std_logic_vector(33 downto 0) := (others => '0');
signal s718 : std_logic_vector(33 downto 0) := (others => '0');
signal s719 : std_logic_vector(33 downto 0) := (others => '0');
signal s720 : std_logic_vector(33 downto 0) := (others => '0');
signal s721 : std_logic_vector(33 downto 0) := (others => '0');
signal s722 : std_logic_vector(33 downto 0) := (others => '0');
signal s723 : std_logic_vector(33 downto 0) := (others => '0');
signal s724 : std_logic_vector(33 downto 0) := (others => '0');
signal s725 : std_logic_vector(33 downto 0) := (others => '0');
signal s726 : std_logic_vector(33 downto 0) := (others => '0');
signal s727 : std_logic_vector(33 downto 0) := (others => '0');
signal s728 : std_logic_vector(33 downto 0) := (others => '0');
signal s729 : std_logic_vector(33 downto 0) := (others => '0');
signal s730 : std_logic_vector(33 downto 0) := (others => '0');
signal s731 : std_logic_vector(33 downto 0) := (others => '0');
signal s732 : std_logic_vector(33 downto 0) := (others => '0');
signal s733 : std_logic_vector(33 downto 0) := (others => '0');
signal s734 : std_logic_vector(33 downto 0) := (others => '0');
signal s735 : std_logic_vector(33 downto 0) := (others => '0');
signal s736 : std_logic_vector(33 downto 0) := (others => '0');
signal s737 : std_logic_vector(33 downto 0) := (others => '0');
signal s738 : std_logic_vector(33 downto 0) := (others => '0');
signal s739 : std_logic_vector(33 downto 0) := (others => '0');
signal s740 : std_logic_vector(33 downto 0) := (others => '0');
signal s741 : std_logic_vector(33 downto 0) := (others => '0');
signal s742 : std_logic_vector(33 downto 0) := (others => '0');
signal s743 : std_logic_vector(33 downto 0) := (others => '0');
signal s744 : std_logic_vector(33 downto 0) := (others => '0');
signal s745 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
      s558 <= "0000000000000000000000000000000000";
      s559 <= "0000000000000000000000000000000000";
      s560 <= "0000000000000000000000000000000000";
      s561 <= "0000000000000000000000000000000000";
      s562 <= "0000000000000000000000000000000000";
      s563 <= "0000000000000000000000000000000000";
      s564 <= "0000000000000000000000000000000000";
      s565 <= "0000000000000000000000000000000000";
      s566 <= "0000000000000000000000000000000000";
      s567 <= "0000000000000000000000000000000000";
      s568 <= "0000000000000000000000000000000000";
      s569 <= "0000000000000000000000000000000000";
      s570 <= "0000000000000000000000000000000000";
      s571 <= "0000000000000000000000000000000000";
      s572 <= "0000000000000000000000000000000000";
      s573 <= "0000000000000000000000000000000000";
      s574 <= "0000000000000000000000000000000000";
      s575 <= "0000000000000000000000000000000000";
      s576 <= "0000000000000000000000000000000000";
      s577 <= "0000000000000000000000000000000000";
      s578 <= "0000000000000000000000000000000000";
      s579 <= "0000000000000000000000000000000000";
      s580 <= "0000000000000000000000000000000000";
      s581 <= "0000000000000000000000000000000000";
      s582 <= "0000000000000000000000000000000000";
      s583 <= "0000000000000000000000000000000000";
      s584 <= "0000000000000000000000000000000000";
      s585 <= "0000000000000000000000000000000000";
      s586 <= "0000000000000000000000000000000000";
      s587 <= "0000000000000000000000000000000000";
      s588 <= "0000000000000000000000000000000000";
      s589 <= "0000000000000000000000000000000000";
      s590 <= "0000000000000000000000000000000000";
      s591 <= "0000000000000000000000000000000000";
      s592 <= "0000000000000000000000000000000000";
      s593 <= "0000000000000000000000000000000000";
      s594 <= "0000000000000000000000000000000000";
      s595 <= "0000000000000000000000000000000000";
      s596 <= "0000000000000000000000000000000000";
      s597 <= "0000000000000000000000000000000000";
      s598 <= "0000000000000000000000000000000000";
      s599 <= "0000000000000000000000000000000000";
      s600 <= "0000000000000000000000000000000000";
      s601 <= "0000000000000000000000000000000000";
      s602 <= "0000000000000000000000000000000000";
      s603 <= "0000000000000000000000000000000000";
      s604 <= "0000000000000000000000000000000000";
      s605 <= "0000000000000000000000000000000000";
      s606 <= "0000000000000000000000000000000000";
      s607 <= "0000000000000000000000000000000000";
      s608 <= "0000000000000000000000000000000000";
      s609 <= "0000000000000000000000000000000000";
      s610 <= "0000000000000000000000000000000000";
      s611 <= "0000000000000000000000000000000000";
      s612 <= "0000000000000000000000000000000000";
      s613 <= "0000000000000000000000000000000000";
      s614 <= "0000000000000000000000000000000000";
      s615 <= "0000000000000000000000000000000000";
      s616 <= "0000000000000000000000000000000000";
      s617 <= "0000000000000000000000000000000000";
      s618 <= "0000000000000000000000000000000000";
      s619 <= "0000000000000000000000000000000000";
      s620 <= "0000000000000000000000000000000000";
      s621 <= "0000000000000000000000000000000000";
      s622 <= "0000000000000000000000000000000000";
      s623 <= "0000000000000000000000000000000000";
      s624 <= "0000000000000000000000000000000000";
      s625 <= "0000000000000000000000000000000000";
      s626 <= "0000000000000000000000000000000000";
      s627 <= "0000000000000000000000000000000000";
      s628 <= "0000000000000000000000000000000000";
      s629 <= "0000000000000000000000000000000000";
      s630 <= "0000000000000000000000000000000000";
      s631 <= "0000000000000000000000000000000000";
      s632 <= "0000000000000000000000000000000000";
      s633 <= "0000000000000000000000000000000000";
      s634 <= "0000000000000000000000000000000000";
      s635 <= "0000000000000000000000000000000000";
      s636 <= "0000000000000000000000000000000000";
      s637 <= "0000000000000000000000000000000000";
      s638 <= "0000000000000000000000000000000000";
      s639 <= "0000000000000000000000000000000000";
      s640 <= "0000000000000000000000000000000000";
      s641 <= "0000000000000000000000000000000000";
      s642 <= "0000000000000000000000000000000000";
      s643 <= "0000000000000000000000000000000000";
      s644 <= "0000000000000000000000000000000000";
      s645 <= "0000000000000000000000000000000000";
      s646 <= "0000000000000000000000000000000000";
      s647 <= "0000000000000000000000000000000000";
      s648 <= "0000000000000000000000000000000000";
      s649 <= "0000000000000000000000000000000000";
      s650 <= "0000000000000000000000000000000000";
      s651 <= "0000000000000000000000000000000000";
      s652 <= "0000000000000000000000000000000000";
      s653 <= "0000000000000000000000000000000000";
      s654 <= "0000000000000000000000000000000000";
      s655 <= "0000000000000000000000000000000000";
      s656 <= "0000000000000000000000000000000000";
      s657 <= "0000000000000000000000000000000000";
      s658 <= "0000000000000000000000000000000000";
      s659 <= "0000000000000000000000000000000000";
      s660 <= "0000000000000000000000000000000000";
      s661 <= "0000000000000000000000000000000000";
      s662 <= "0000000000000000000000000000000000";
      s663 <= "0000000000000000000000000000000000";
      s664 <= "0000000000000000000000000000000000";
      s665 <= "0000000000000000000000000000000000";
      s666 <= "0000000000000000000000000000000000";
      s667 <= "0000000000000000000000000000000000";
      s668 <= "0000000000000000000000000000000000";
      s669 <= "0000000000000000000000000000000000";
      s670 <= "0000000000000000000000000000000000";
      s671 <= "0000000000000000000000000000000000";
      s672 <= "0000000000000000000000000000000000";
      s673 <= "0000000000000000000000000000000000";
      s674 <= "0000000000000000000000000000000000";
      s675 <= "0000000000000000000000000000000000";
      s676 <= "0000000000000000000000000000000000";
      s677 <= "0000000000000000000000000000000000";
      s678 <= "0000000000000000000000000000000000";
      s679 <= "0000000000000000000000000000000000";
      s680 <= "0000000000000000000000000000000000";
      s681 <= "0000000000000000000000000000000000";
      s682 <= "0000000000000000000000000000000000";
      s683 <= "0000000000000000000000000000000000";
      s684 <= "0000000000000000000000000000000000";
      s685 <= "0000000000000000000000000000000000";
      s686 <= "0000000000000000000000000000000000";
      s687 <= "0000000000000000000000000000000000";
      s688 <= "0000000000000000000000000000000000";
      s689 <= "0000000000000000000000000000000000";
      s690 <= "0000000000000000000000000000000000";
      s691 <= "0000000000000000000000000000000000";
      s692 <= "0000000000000000000000000000000000";
      s693 <= "0000000000000000000000000000000000";
      s694 <= "0000000000000000000000000000000000";
      s695 <= "0000000000000000000000000000000000";
      s696 <= "0000000000000000000000000000000000";
      s697 <= "0000000000000000000000000000000000";
      s698 <= "0000000000000000000000000000000000";
      s699 <= "0000000000000000000000000000000000";
      s700 <= "0000000000000000000000000000000000";
      s701 <= "0000000000000000000000000000000000";
      s702 <= "0000000000000000000000000000000000";
      s703 <= "0000000000000000000000000000000000";
      s704 <= "0000000000000000000000000000000000";
      s705 <= "0000000000000000000000000000000000";
      s706 <= "0000000000000000000000000000000000";
      s707 <= "0000000000000000000000000000000000";
      s708 <= "0000000000000000000000000000000000";
      s709 <= "0000000000000000000000000000000000";
      s710 <= "0000000000000000000000000000000000";
      s711 <= "0000000000000000000000000000000000";
      s712 <= "0000000000000000000000000000000000";
      s713 <= "0000000000000000000000000000000000";
      s714 <= "0000000000000000000000000000000000";
      s715 <= "0000000000000000000000000000000000";
      s716 <= "0000000000000000000000000000000000";
      s717 <= "0000000000000000000000000000000000";
      s718 <= "0000000000000000000000000000000000";
      s719 <= "0000000000000000000000000000000000";
      s720 <= "0000000000000000000000000000000000";
      s721 <= "0000000000000000000000000000000000";
      s722 <= "0000000000000000000000000000000000";
      s723 <= "0000000000000000000000000000000000";
      s724 <= "0000000000000000000000000000000000";
      s725 <= "0000000000000000000000000000000000";
      s726 <= "0000000000000000000000000000000000";
      s727 <= "0000000000000000000000000000000000";
      s728 <= "0000000000000000000000000000000000";
      s729 <= "0000000000000000000000000000000000";
      s730 <= "0000000000000000000000000000000000";
      s731 <= "0000000000000000000000000000000000";
      s732 <= "0000000000000000000000000000000000";
      s733 <= "0000000000000000000000000000000000";
      s734 <= "0000000000000000000000000000000000";
      s735 <= "0000000000000000000000000000000000";
      s736 <= "0000000000000000000000000000000000";
      s737 <= "0000000000000000000000000000000000";
      s738 <= "0000000000000000000000000000000000";
      s739 <= "0000000000000000000000000000000000";
      s740 <= "0000000000000000000000000000000000";
      s741 <= "0000000000000000000000000000000000";
      s742 <= "0000000000000000000000000000000000";
      s743 <= "0000000000000000000000000000000000";
      s744 <= "0000000000000000000000000000000000";
      s745 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      s558 <= s557;
      s559 <= s558;
      s560 <= s559;
      s561 <= s560;
      s562 <= s561;
      s563 <= s562;
      s564 <= s563;
      s565 <= s564;
      s566 <= s565;
      s567 <= s566;
      s568 <= s567;
      s569 <= s568;
      s570 <= s569;
      s571 <= s570;
      s572 <= s571;
      s573 <= s572;
      s574 <= s573;
      s575 <= s574;
      s576 <= s575;
      s577 <= s576;
      s578 <= s577;
      s579 <= s578;
      s580 <= s579;
      s581 <= s580;
      s582 <= s581;
      s583 <= s582;
      s584 <= s583;
      s585 <= s584;
      s586 <= s585;
      s587 <= s586;
      s588 <= s587;
      s589 <= s588;
      s590 <= s589;
      s591 <= s590;
      s592 <= s591;
      s593 <= s592;
      s594 <= s593;
      s595 <= s594;
      s596 <= s595;
      s597 <= s596;
      s598 <= s597;
      s599 <= s598;
      s600 <= s599;
      s601 <= s600;
      s602 <= s601;
      s603 <= s602;
      s604 <= s603;
      s605 <= s604;
      s606 <= s605;
      s607 <= s606;
      s608 <= s607;
      s609 <= s608;
      s610 <= s609;
      s611 <= s610;
      s612 <= s611;
      s613 <= s612;
      s614 <= s613;
      s615 <= s614;
      s616 <= s615;
      s617 <= s616;
      s618 <= s617;
      s619 <= s618;
      s620 <= s619;
      s621 <= s620;
      s622 <= s621;
      s623 <= s622;
      s624 <= s623;
      s625 <= s624;
      s626 <= s625;
      s627 <= s626;
      s628 <= s627;
      s629 <= s628;
      s630 <= s629;
      s631 <= s630;
      s632 <= s631;
      s633 <= s632;
      s634 <= s633;
      s635 <= s634;
      s636 <= s635;
      s637 <= s636;
      s638 <= s637;
      s639 <= s638;
      s640 <= s639;
      s641 <= s640;
      s642 <= s641;
      s643 <= s642;
      s644 <= s643;
      s645 <= s644;
      s646 <= s645;
      s647 <= s646;
      s648 <= s647;
      s649 <= s648;
      s650 <= s649;
      s651 <= s650;
      s652 <= s651;
      s653 <= s652;
      s654 <= s653;
      s655 <= s654;
      s656 <= s655;
      s657 <= s656;
      s658 <= s657;
      s659 <= s658;
      s660 <= s659;
      s661 <= s660;
      s662 <= s661;
      s663 <= s662;
      s664 <= s663;
      s665 <= s664;
      s666 <= s665;
      s667 <= s666;
      s668 <= s667;
      s669 <= s668;
      s670 <= s669;
      s671 <= s670;
      s672 <= s671;
      s673 <= s672;
      s674 <= s673;
      s675 <= s674;
      s676 <= s675;
      s677 <= s676;
      s678 <= s677;
      s679 <= s678;
      s680 <= s679;
      s681 <= s680;
      s682 <= s681;
      s683 <= s682;
      s684 <= s683;
      s685 <= s684;
      s686 <= s685;
      s687 <= s686;
      s688 <= s687;
      s689 <= s688;
      s690 <= s689;
      s691 <= s690;
      s692 <= s691;
      s693 <= s692;
      s694 <= s693;
      s695 <= s694;
      s696 <= s695;
      s697 <= s696;
      s698 <= s697;
      s699 <= s698;
      s700 <= s699;
      s701 <= s700;
      s702 <= s701;
      s703 <= s702;
      s704 <= s703;
      s705 <= s704;
      s706 <= s705;
      s707 <= s706;
      s708 <= s707;
      s709 <= s708;
      s710 <= s709;
      s711 <= s710;
      s712 <= s711;
      s713 <= s712;
      s714 <= s713;
      s715 <= s714;
      s716 <= s715;
      s717 <= s716;
      s718 <= s717;
      s719 <= s718;
      s720 <= s719;
      s721 <= s720;
      s722 <= s721;
      s723 <= s722;
      s724 <= s723;
      s725 <= s724;
      s726 <= s725;
      s727 <= s726;
      s728 <= s727;
      s729 <= s728;
      s730 <= s729;
      s731 <= s730;
      s732 <= s731;
      s733 <= s732;
      s734 <= s733;
      s735 <= s734;
      s736 <= s735;
      s737 <= s736;
      s738 <= s737;
      s739 <= s738;
      s740 <= s739;
      s741 <= s740;
      s742 <= s741;
      s743 <= s742;
      s744 <= s743;
      s745 <= s744;
      Y <= s745;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_849_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 849 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_849_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_849_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
signal s558 : std_logic_vector(33 downto 0) := (others => '0');
signal s559 : std_logic_vector(33 downto 0) := (others => '0');
signal s560 : std_logic_vector(33 downto 0) := (others => '0');
signal s561 : std_logic_vector(33 downto 0) := (others => '0');
signal s562 : std_logic_vector(33 downto 0) := (others => '0');
signal s563 : std_logic_vector(33 downto 0) := (others => '0');
signal s564 : std_logic_vector(33 downto 0) := (others => '0');
signal s565 : std_logic_vector(33 downto 0) := (others => '0');
signal s566 : std_logic_vector(33 downto 0) := (others => '0');
signal s567 : std_logic_vector(33 downto 0) := (others => '0');
signal s568 : std_logic_vector(33 downto 0) := (others => '0');
signal s569 : std_logic_vector(33 downto 0) := (others => '0');
signal s570 : std_logic_vector(33 downto 0) := (others => '0');
signal s571 : std_logic_vector(33 downto 0) := (others => '0');
signal s572 : std_logic_vector(33 downto 0) := (others => '0');
signal s573 : std_logic_vector(33 downto 0) := (others => '0');
signal s574 : std_logic_vector(33 downto 0) := (others => '0');
signal s575 : std_logic_vector(33 downto 0) := (others => '0');
signal s576 : std_logic_vector(33 downto 0) := (others => '0');
signal s577 : std_logic_vector(33 downto 0) := (others => '0');
signal s578 : std_logic_vector(33 downto 0) := (others => '0');
signal s579 : std_logic_vector(33 downto 0) := (others => '0');
signal s580 : std_logic_vector(33 downto 0) := (others => '0');
signal s581 : std_logic_vector(33 downto 0) := (others => '0');
signal s582 : std_logic_vector(33 downto 0) := (others => '0');
signal s583 : std_logic_vector(33 downto 0) := (others => '0');
signal s584 : std_logic_vector(33 downto 0) := (others => '0');
signal s585 : std_logic_vector(33 downto 0) := (others => '0');
signal s586 : std_logic_vector(33 downto 0) := (others => '0');
signal s587 : std_logic_vector(33 downto 0) := (others => '0');
signal s588 : std_logic_vector(33 downto 0) := (others => '0');
signal s589 : std_logic_vector(33 downto 0) := (others => '0');
signal s590 : std_logic_vector(33 downto 0) := (others => '0');
signal s591 : std_logic_vector(33 downto 0) := (others => '0');
signal s592 : std_logic_vector(33 downto 0) := (others => '0');
signal s593 : std_logic_vector(33 downto 0) := (others => '0');
signal s594 : std_logic_vector(33 downto 0) := (others => '0');
signal s595 : std_logic_vector(33 downto 0) := (others => '0');
signal s596 : std_logic_vector(33 downto 0) := (others => '0');
signal s597 : std_logic_vector(33 downto 0) := (others => '0');
signal s598 : std_logic_vector(33 downto 0) := (others => '0');
signal s599 : std_logic_vector(33 downto 0) := (others => '0');
signal s600 : std_logic_vector(33 downto 0) := (others => '0');
signal s601 : std_logic_vector(33 downto 0) := (others => '0');
signal s602 : std_logic_vector(33 downto 0) := (others => '0');
signal s603 : std_logic_vector(33 downto 0) := (others => '0');
signal s604 : std_logic_vector(33 downto 0) := (others => '0');
signal s605 : std_logic_vector(33 downto 0) := (others => '0');
signal s606 : std_logic_vector(33 downto 0) := (others => '0');
signal s607 : std_logic_vector(33 downto 0) := (others => '0');
signal s608 : std_logic_vector(33 downto 0) := (others => '0');
signal s609 : std_logic_vector(33 downto 0) := (others => '0');
signal s610 : std_logic_vector(33 downto 0) := (others => '0');
signal s611 : std_logic_vector(33 downto 0) := (others => '0');
signal s612 : std_logic_vector(33 downto 0) := (others => '0');
signal s613 : std_logic_vector(33 downto 0) := (others => '0');
signal s614 : std_logic_vector(33 downto 0) := (others => '0');
signal s615 : std_logic_vector(33 downto 0) := (others => '0');
signal s616 : std_logic_vector(33 downto 0) := (others => '0');
signal s617 : std_logic_vector(33 downto 0) := (others => '0');
signal s618 : std_logic_vector(33 downto 0) := (others => '0');
signal s619 : std_logic_vector(33 downto 0) := (others => '0');
signal s620 : std_logic_vector(33 downto 0) := (others => '0');
signal s621 : std_logic_vector(33 downto 0) := (others => '0');
signal s622 : std_logic_vector(33 downto 0) := (others => '0');
signal s623 : std_logic_vector(33 downto 0) := (others => '0');
signal s624 : std_logic_vector(33 downto 0) := (others => '0');
signal s625 : std_logic_vector(33 downto 0) := (others => '0');
signal s626 : std_logic_vector(33 downto 0) := (others => '0');
signal s627 : std_logic_vector(33 downto 0) := (others => '0');
signal s628 : std_logic_vector(33 downto 0) := (others => '0');
signal s629 : std_logic_vector(33 downto 0) := (others => '0');
signal s630 : std_logic_vector(33 downto 0) := (others => '0');
signal s631 : std_logic_vector(33 downto 0) := (others => '0');
signal s632 : std_logic_vector(33 downto 0) := (others => '0');
signal s633 : std_logic_vector(33 downto 0) := (others => '0');
signal s634 : std_logic_vector(33 downto 0) := (others => '0');
signal s635 : std_logic_vector(33 downto 0) := (others => '0');
signal s636 : std_logic_vector(33 downto 0) := (others => '0');
signal s637 : std_logic_vector(33 downto 0) := (others => '0');
signal s638 : std_logic_vector(33 downto 0) := (others => '0');
signal s639 : std_logic_vector(33 downto 0) := (others => '0');
signal s640 : std_logic_vector(33 downto 0) := (others => '0');
signal s641 : std_logic_vector(33 downto 0) := (others => '0');
signal s642 : std_logic_vector(33 downto 0) := (others => '0');
signal s643 : std_logic_vector(33 downto 0) := (others => '0');
signal s644 : std_logic_vector(33 downto 0) := (others => '0');
signal s645 : std_logic_vector(33 downto 0) := (others => '0');
signal s646 : std_logic_vector(33 downto 0) := (others => '0');
signal s647 : std_logic_vector(33 downto 0) := (others => '0');
signal s648 : std_logic_vector(33 downto 0) := (others => '0');
signal s649 : std_logic_vector(33 downto 0) := (others => '0');
signal s650 : std_logic_vector(33 downto 0) := (others => '0');
signal s651 : std_logic_vector(33 downto 0) := (others => '0');
signal s652 : std_logic_vector(33 downto 0) := (others => '0');
signal s653 : std_logic_vector(33 downto 0) := (others => '0');
signal s654 : std_logic_vector(33 downto 0) := (others => '0');
signal s655 : std_logic_vector(33 downto 0) := (others => '0');
signal s656 : std_logic_vector(33 downto 0) := (others => '0');
signal s657 : std_logic_vector(33 downto 0) := (others => '0');
signal s658 : std_logic_vector(33 downto 0) := (others => '0');
signal s659 : std_logic_vector(33 downto 0) := (others => '0');
signal s660 : std_logic_vector(33 downto 0) := (others => '0');
signal s661 : std_logic_vector(33 downto 0) := (others => '0');
signal s662 : std_logic_vector(33 downto 0) := (others => '0');
signal s663 : std_logic_vector(33 downto 0) := (others => '0');
signal s664 : std_logic_vector(33 downto 0) := (others => '0');
signal s665 : std_logic_vector(33 downto 0) := (others => '0');
signal s666 : std_logic_vector(33 downto 0) := (others => '0');
signal s667 : std_logic_vector(33 downto 0) := (others => '0');
signal s668 : std_logic_vector(33 downto 0) := (others => '0');
signal s669 : std_logic_vector(33 downto 0) := (others => '0');
signal s670 : std_logic_vector(33 downto 0) := (others => '0');
signal s671 : std_logic_vector(33 downto 0) := (others => '0');
signal s672 : std_logic_vector(33 downto 0) := (others => '0');
signal s673 : std_logic_vector(33 downto 0) := (others => '0');
signal s674 : std_logic_vector(33 downto 0) := (others => '0');
signal s675 : std_logic_vector(33 downto 0) := (others => '0');
signal s676 : std_logic_vector(33 downto 0) := (others => '0');
signal s677 : std_logic_vector(33 downto 0) := (others => '0');
signal s678 : std_logic_vector(33 downto 0) := (others => '0');
signal s679 : std_logic_vector(33 downto 0) := (others => '0');
signal s680 : std_logic_vector(33 downto 0) := (others => '0');
signal s681 : std_logic_vector(33 downto 0) := (others => '0');
signal s682 : std_logic_vector(33 downto 0) := (others => '0');
signal s683 : std_logic_vector(33 downto 0) := (others => '0');
signal s684 : std_logic_vector(33 downto 0) := (others => '0');
signal s685 : std_logic_vector(33 downto 0) := (others => '0');
signal s686 : std_logic_vector(33 downto 0) := (others => '0');
signal s687 : std_logic_vector(33 downto 0) := (others => '0');
signal s688 : std_logic_vector(33 downto 0) := (others => '0');
signal s689 : std_logic_vector(33 downto 0) := (others => '0');
signal s690 : std_logic_vector(33 downto 0) := (others => '0');
signal s691 : std_logic_vector(33 downto 0) := (others => '0');
signal s692 : std_logic_vector(33 downto 0) := (others => '0');
signal s693 : std_logic_vector(33 downto 0) := (others => '0');
signal s694 : std_logic_vector(33 downto 0) := (others => '0');
signal s695 : std_logic_vector(33 downto 0) := (others => '0');
signal s696 : std_logic_vector(33 downto 0) := (others => '0');
signal s697 : std_logic_vector(33 downto 0) := (others => '0');
signal s698 : std_logic_vector(33 downto 0) := (others => '0');
signal s699 : std_logic_vector(33 downto 0) := (others => '0');
signal s700 : std_logic_vector(33 downto 0) := (others => '0');
signal s701 : std_logic_vector(33 downto 0) := (others => '0');
signal s702 : std_logic_vector(33 downto 0) := (others => '0');
signal s703 : std_logic_vector(33 downto 0) := (others => '0');
signal s704 : std_logic_vector(33 downto 0) := (others => '0');
signal s705 : std_logic_vector(33 downto 0) := (others => '0');
signal s706 : std_logic_vector(33 downto 0) := (others => '0');
signal s707 : std_logic_vector(33 downto 0) := (others => '0');
signal s708 : std_logic_vector(33 downto 0) := (others => '0');
signal s709 : std_logic_vector(33 downto 0) := (others => '0');
signal s710 : std_logic_vector(33 downto 0) := (others => '0');
signal s711 : std_logic_vector(33 downto 0) := (others => '0');
signal s712 : std_logic_vector(33 downto 0) := (others => '0');
signal s713 : std_logic_vector(33 downto 0) := (others => '0');
signal s714 : std_logic_vector(33 downto 0) := (others => '0');
signal s715 : std_logic_vector(33 downto 0) := (others => '0');
signal s716 : std_logic_vector(33 downto 0) := (others => '0');
signal s717 : std_logic_vector(33 downto 0) := (others => '0');
signal s718 : std_logic_vector(33 downto 0) := (others => '0');
signal s719 : std_logic_vector(33 downto 0) := (others => '0');
signal s720 : std_logic_vector(33 downto 0) := (others => '0');
signal s721 : std_logic_vector(33 downto 0) := (others => '0');
signal s722 : std_logic_vector(33 downto 0) := (others => '0');
signal s723 : std_logic_vector(33 downto 0) := (others => '0');
signal s724 : std_logic_vector(33 downto 0) := (others => '0');
signal s725 : std_logic_vector(33 downto 0) := (others => '0');
signal s726 : std_logic_vector(33 downto 0) := (others => '0');
signal s727 : std_logic_vector(33 downto 0) := (others => '0');
signal s728 : std_logic_vector(33 downto 0) := (others => '0');
signal s729 : std_logic_vector(33 downto 0) := (others => '0');
signal s730 : std_logic_vector(33 downto 0) := (others => '0');
signal s731 : std_logic_vector(33 downto 0) := (others => '0');
signal s732 : std_logic_vector(33 downto 0) := (others => '0');
signal s733 : std_logic_vector(33 downto 0) := (others => '0');
signal s734 : std_logic_vector(33 downto 0) := (others => '0');
signal s735 : std_logic_vector(33 downto 0) := (others => '0');
signal s736 : std_logic_vector(33 downto 0) := (others => '0');
signal s737 : std_logic_vector(33 downto 0) := (others => '0');
signal s738 : std_logic_vector(33 downto 0) := (others => '0');
signal s739 : std_logic_vector(33 downto 0) := (others => '0');
signal s740 : std_logic_vector(33 downto 0) := (others => '0');
signal s741 : std_logic_vector(33 downto 0) := (others => '0');
signal s742 : std_logic_vector(33 downto 0) := (others => '0');
signal s743 : std_logic_vector(33 downto 0) := (others => '0');
signal s744 : std_logic_vector(33 downto 0) := (others => '0');
signal s745 : std_logic_vector(33 downto 0) := (others => '0');
signal s746 : std_logic_vector(33 downto 0) := (others => '0');
signal s747 : std_logic_vector(33 downto 0) := (others => '0');
signal s748 : std_logic_vector(33 downto 0) := (others => '0');
signal s749 : std_logic_vector(33 downto 0) := (others => '0');
signal s750 : std_logic_vector(33 downto 0) := (others => '0');
signal s751 : std_logic_vector(33 downto 0) := (others => '0');
signal s752 : std_logic_vector(33 downto 0) := (others => '0');
signal s753 : std_logic_vector(33 downto 0) := (others => '0');
signal s754 : std_logic_vector(33 downto 0) := (others => '0');
signal s755 : std_logic_vector(33 downto 0) := (others => '0');
signal s756 : std_logic_vector(33 downto 0) := (others => '0');
signal s757 : std_logic_vector(33 downto 0) := (others => '0');
signal s758 : std_logic_vector(33 downto 0) := (others => '0');
signal s759 : std_logic_vector(33 downto 0) := (others => '0');
signal s760 : std_logic_vector(33 downto 0) := (others => '0');
signal s761 : std_logic_vector(33 downto 0) := (others => '0');
signal s762 : std_logic_vector(33 downto 0) := (others => '0');
signal s763 : std_logic_vector(33 downto 0) := (others => '0');
signal s764 : std_logic_vector(33 downto 0) := (others => '0');
signal s765 : std_logic_vector(33 downto 0) := (others => '0');
signal s766 : std_logic_vector(33 downto 0) := (others => '0');
signal s767 : std_logic_vector(33 downto 0) := (others => '0');
signal s768 : std_logic_vector(33 downto 0) := (others => '0');
signal s769 : std_logic_vector(33 downto 0) := (others => '0');
signal s770 : std_logic_vector(33 downto 0) := (others => '0');
signal s771 : std_logic_vector(33 downto 0) := (others => '0');
signal s772 : std_logic_vector(33 downto 0) := (others => '0');
signal s773 : std_logic_vector(33 downto 0) := (others => '0');
signal s774 : std_logic_vector(33 downto 0) := (others => '0');
signal s775 : std_logic_vector(33 downto 0) := (others => '0');
signal s776 : std_logic_vector(33 downto 0) := (others => '0');
signal s777 : std_logic_vector(33 downto 0) := (others => '0');
signal s778 : std_logic_vector(33 downto 0) := (others => '0');
signal s779 : std_logic_vector(33 downto 0) := (others => '0');
signal s780 : std_logic_vector(33 downto 0) := (others => '0');
signal s781 : std_logic_vector(33 downto 0) := (others => '0');
signal s782 : std_logic_vector(33 downto 0) := (others => '0');
signal s783 : std_logic_vector(33 downto 0) := (others => '0');
signal s784 : std_logic_vector(33 downto 0) := (others => '0');
signal s785 : std_logic_vector(33 downto 0) := (others => '0');
signal s786 : std_logic_vector(33 downto 0) := (others => '0');
signal s787 : std_logic_vector(33 downto 0) := (others => '0');
signal s788 : std_logic_vector(33 downto 0) := (others => '0');
signal s789 : std_logic_vector(33 downto 0) := (others => '0');
signal s790 : std_logic_vector(33 downto 0) := (others => '0');
signal s791 : std_logic_vector(33 downto 0) := (others => '0');
signal s792 : std_logic_vector(33 downto 0) := (others => '0');
signal s793 : std_logic_vector(33 downto 0) := (others => '0');
signal s794 : std_logic_vector(33 downto 0) := (others => '0');
signal s795 : std_logic_vector(33 downto 0) := (others => '0');
signal s796 : std_logic_vector(33 downto 0) := (others => '0');
signal s797 : std_logic_vector(33 downto 0) := (others => '0');
signal s798 : std_logic_vector(33 downto 0) := (others => '0');
signal s799 : std_logic_vector(33 downto 0) := (others => '0');
signal s800 : std_logic_vector(33 downto 0) := (others => '0');
signal s801 : std_logic_vector(33 downto 0) := (others => '0');
signal s802 : std_logic_vector(33 downto 0) := (others => '0');
signal s803 : std_logic_vector(33 downto 0) := (others => '0');
signal s804 : std_logic_vector(33 downto 0) := (others => '0');
signal s805 : std_logic_vector(33 downto 0) := (others => '0');
signal s806 : std_logic_vector(33 downto 0) := (others => '0');
signal s807 : std_logic_vector(33 downto 0) := (others => '0');
signal s808 : std_logic_vector(33 downto 0) := (others => '0');
signal s809 : std_logic_vector(33 downto 0) := (others => '0');
signal s810 : std_logic_vector(33 downto 0) := (others => '0');
signal s811 : std_logic_vector(33 downto 0) := (others => '0');
signal s812 : std_logic_vector(33 downto 0) := (others => '0');
signal s813 : std_logic_vector(33 downto 0) := (others => '0');
signal s814 : std_logic_vector(33 downto 0) := (others => '0');
signal s815 : std_logic_vector(33 downto 0) := (others => '0');
signal s816 : std_logic_vector(33 downto 0) := (others => '0');
signal s817 : std_logic_vector(33 downto 0) := (others => '0');
signal s818 : std_logic_vector(33 downto 0) := (others => '0');
signal s819 : std_logic_vector(33 downto 0) := (others => '0');
signal s820 : std_logic_vector(33 downto 0) := (others => '0');
signal s821 : std_logic_vector(33 downto 0) := (others => '0');
signal s822 : std_logic_vector(33 downto 0) := (others => '0');
signal s823 : std_logic_vector(33 downto 0) := (others => '0');
signal s824 : std_logic_vector(33 downto 0) := (others => '0');
signal s825 : std_logic_vector(33 downto 0) := (others => '0');
signal s826 : std_logic_vector(33 downto 0) := (others => '0');
signal s827 : std_logic_vector(33 downto 0) := (others => '0');
signal s828 : std_logic_vector(33 downto 0) := (others => '0');
signal s829 : std_logic_vector(33 downto 0) := (others => '0');
signal s830 : std_logic_vector(33 downto 0) := (others => '0');
signal s831 : std_logic_vector(33 downto 0) := (others => '0');
signal s832 : std_logic_vector(33 downto 0) := (others => '0');
signal s833 : std_logic_vector(33 downto 0) := (others => '0');
signal s834 : std_logic_vector(33 downto 0) := (others => '0');
signal s835 : std_logic_vector(33 downto 0) := (others => '0');
signal s836 : std_logic_vector(33 downto 0) := (others => '0');
signal s837 : std_logic_vector(33 downto 0) := (others => '0');
signal s838 : std_logic_vector(33 downto 0) := (others => '0');
signal s839 : std_logic_vector(33 downto 0) := (others => '0');
signal s840 : std_logic_vector(33 downto 0) := (others => '0');
signal s841 : std_logic_vector(33 downto 0) := (others => '0');
signal s842 : std_logic_vector(33 downto 0) := (others => '0');
signal s843 : std_logic_vector(33 downto 0) := (others => '0');
signal s844 : std_logic_vector(33 downto 0) := (others => '0');
signal s845 : std_logic_vector(33 downto 0) := (others => '0');
signal s846 : std_logic_vector(33 downto 0) := (others => '0');
signal s847 : std_logic_vector(33 downto 0) := (others => '0');
signal s848 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
      s558 <= "0000000000000000000000000000000000";
      s559 <= "0000000000000000000000000000000000";
      s560 <= "0000000000000000000000000000000000";
      s561 <= "0000000000000000000000000000000000";
      s562 <= "0000000000000000000000000000000000";
      s563 <= "0000000000000000000000000000000000";
      s564 <= "0000000000000000000000000000000000";
      s565 <= "0000000000000000000000000000000000";
      s566 <= "0000000000000000000000000000000000";
      s567 <= "0000000000000000000000000000000000";
      s568 <= "0000000000000000000000000000000000";
      s569 <= "0000000000000000000000000000000000";
      s570 <= "0000000000000000000000000000000000";
      s571 <= "0000000000000000000000000000000000";
      s572 <= "0000000000000000000000000000000000";
      s573 <= "0000000000000000000000000000000000";
      s574 <= "0000000000000000000000000000000000";
      s575 <= "0000000000000000000000000000000000";
      s576 <= "0000000000000000000000000000000000";
      s577 <= "0000000000000000000000000000000000";
      s578 <= "0000000000000000000000000000000000";
      s579 <= "0000000000000000000000000000000000";
      s580 <= "0000000000000000000000000000000000";
      s581 <= "0000000000000000000000000000000000";
      s582 <= "0000000000000000000000000000000000";
      s583 <= "0000000000000000000000000000000000";
      s584 <= "0000000000000000000000000000000000";
      s585 <= "0000000000000000000000000000000000";
      s586 <= "0000000000000000000000000000000000";
      s587 <= "0000000000000000000000000000000000";
      s588 <= "0000000000000000000000000000000000";
      s589 <= "0000000000000000000000000000000000";
      s590 <= "0000000000000000000000000000000000";
      s591 <= "0000000000000000000000000000000000";
      s592 <= "0000000000000000000000000000000000";
      s593 <= "0000000000000000000000000000000000";
      s594 <= "0000000000000000000000000000000000";
      s595 <= "0000000000000000000000000000000000";
      s596 <= "0000000000000000000000000000000000";
      s597 <= "0000000000000000000000000000000000";
      s598 <= "0000000000000000000000000000000000";
      s599 <= "0000000000000000000000000000000000";
      s600 <= "0000000000000000000000000000000000";
      s601 <= "0000000000000000000000000000000000";
      s602 <= "0000000000000000000000000000000000";
      s603 <= "0000000000000000000000000000000000";
      s604 <= "0000000000000000000000000000000000";
      s605 <= "0000000000000000000000000000000000";
      s606 <= "0000000000000000000000000000000000";
      s607 <= "0000000000000000000000000000000000";
      s608 <= "0000000000000000000000000000000000";
      s609 <= "0000000000000000000000000000000000";
      s610 <= "0000000000000000000000000000000000";
      s611 <= "0000000000000000000000000000000000";
      s612 <= "0000000000000000000000000000000000";
      s613 <= "0000000000000000000000000000000000";
      s614 <= "0000000000000000000000000000000000";
      s615 <= "0000000000000000000000000000000000";
      s616 <= "0000000000000000000000000000000000";
      s617 <= "0000000000000000000000000000000000";
      s618 <= "0000000000000000000000000000000000";
      s619 <= "0000000000000000000000000000000000";
      s620 <= "0000000000000000000000000000000000";
      s621 <= "0000000000000000000000000000000000";
      s622 <= "0000000000000000000000000000000000";
      s623 <= "0000000000000000000000000000000000";
      s624 <= "0000000000000000000000000000000000";
      s625 <= "0000000000000000000000000000000000";
      s626 <= "0000000000000000000000000000000000";
      s627 <= "0000000000000000000000000000000000";
      s628 <= "0000000000000000000000000000000000";
      s629 <= "0000000000000000000000000000000000";
      s630 <= "0000000000000000000000000000000000";
      s631 <= "0000000000000000000000000000000000";
      s632 <= "0000000000000000000000000000000000";
      s633 <= "0000000000000000000000000000000000";
      s634 <= "0000000000000000000000000000000000";
      s635 <= "0000000000000000000000000000000000";
      s636 <= "0000000000000000000000000000000000";
      s637 <= "0000000000000000000000000000000000";
      s638 <= "0000000000000000000000000000000000";
      s639 <= "0000000000000000000000000000000000";
      s640 <= "0000000000000000000000000000000000";
      s641 <= "0000000000000000000000000000000000";
      s642 <= "0000000000000000000000000000000000";
      s643 <= "0000000000000000000000000000000000";
      s644 <= "0000000000000000000000000000000000";
      s645 <= "0000000000000000000000000000000000";
      s646 <= "0000000000000000000000000000000000";
      s647 <= "0000000000000000000000000000000000";
      s648 <= "0000000000000000000000000000000000";
      s649 <= "0000000000000000000000000000000000";
      s650 <= "0000000000000000000000000000000000";
      s651 <= "0000000000000000000000000000000000";
      s652 <= "0000000000000000000000000000000000";
      s653 <= "0000000000000000000000000000000000";
      s654 <= "0000000000000000000000000000000000";
      s655 <= "0000000000000000000000000000000000";
      s656 <= "0000000000000000000000000000000000";
      s657 <= "0000000000000000000000000000000000";
      s658 <= "0000000000000000000000000000000000";
      s659 <= "0000000000000000000000000000000000";
      s660 <= "0000000000000000000000000000000000";
      s661 <= "0000000000000000000000000000000000";
      s662 <= "0000000000000000000000000000000000";
      s663 <= "0000000000000000000000000000000000";
      s664 <= "0000000000000000000000000000000000";
      s665 <= "0000000000000000000000000000000000";
      s666 <= "0000000000000000000000000000000000";
      s667 <= "0000000000000000000000000000000000";
      s668 <= "0000000000000000000000000000000000";
      s669 <= "0000000000000000000000000000000000";
      s670 <= "0000000000000000000000000000000000";
      s671 <= "0000000000000000000000000000000000";
      s672 <= "0000000000000000000000000000000000";
      s673 <= "0000000000000000000000000000000000";
      s674 <= "0000000000000000000000000000000000";
      s675 <= "0000000000000000000000000000000000";
      s676 <= "0000000000000000000000000000000000";
      s677 <= "0000000000000000000000000000000000";
      s678 <= "0000000000000000000000000000000000";
      s679 <= "0000000000000000000000000000000000";
      s680 <= "0000000000000000000000000000000000";
      s681 <= "0000000000000000000000000000000000";
      s682 <= "0000000000000000000000000000000000";
      s683 <= "0000000000000000000000000000000000";
      s684 <= "0000000000000000000000000000000000";
      s685 <= "0000000000000000000000000000000000";
      s686 <= "0000000000000000000000000000000000";
      s687 <= "0000000000000000000000000000000000";
      s688 <= "0000000000000000000000000000000000";
      s689 <= "0000000000000000000000000000000000";
      s690 <= "0000000000000000000000000000000000";
      s691 <= "0000000000000000000000000000000000";
      s692 <= "0000000000000000000000000000000000";
      s693 <= "0000000000000000000000000000000000";
      s694 <= "0000000000000000000000000000000000";
      s695 <= "0000000000000000000000000000000000";
      s696 <= "0000000000000000000000000000000000";
      s697 <= "0000000000000000000000000000000000";
      s698 <= "0000000000000000000000000000000000";
      s699 <= "0000000000000000000000000000000000";
      s700 <= "0000000000000000000000000000000000";
      s701 <= "0000000000000000000000000000000000";
      s702 <= "0000000000000000000000000000000000";
      s703 <= "0000000000000000000000000000000000";
      s704 <= "0000000000000000000000000000000000";
      s705 <= "0000000000000000000000000000000000";
      s706 <= "0000000000000000000000000000000000";
      s707 <= "0000000000000000000000000000000000";
      s708 <= "0000000000000000000000000000000000";
      s709 <= "0000000000000000000000000000000000";
      s710 <= "0000000000000000000000000000000000";
      s711 <= "0000000000000000000000000000000000";
      s712 <= "0000000000000000000000000000000000";
      s713 <= "0000000000000000000000000000000000";
      s714 <= "0000000000000000000000000000000000";
      s715 <= "0000000000000000000000000000000000";
      s716 <= "0000000000000000000000000000000000";
      s717 <= "0000000000000000000000000000000000";
      s718 <= "0000000000000000000000000000000000";
      s719 <= "0000000000000000000000000000000000";
      s720 <= "0000000000000000000000000000000000";
      s721 <= "0000000000000000000000000000000000";
      s722 <= "0000000000000000000000000000000000";
      s723 <= "0000000000000000000000000000000000";
      s724 <= "0000000000000000000000000000000000";
      s725 <= "0000000000000000000000000000000000";
      s726 <= "0000000000000000000000000000000000";
      s727 <= "0000000000000000000000000000000000";
      s728 <= "0000000000000000000000000000000000";
      s729 <= "0000000000000000000000000000000000";
      s730 <= "0000000000000000000000000000000000";
      s731 <= "0000000000000000000000000000000000";
      s732 <= "0000000000000000000000000000000000";
      s733 <= "0000000000000000000000000000000000";
      s734 <= "0000000000000000000000000000000000";
      s735 <= "0000000000000000000000000000000000";
      s736 <= "0000000000000000000000000000000000";
      s737 <= "0000000000000000000000000000000000";
      s738 <= "0000000000000000000000000000000000";
      s739 <= "0000000000000000000000000000000000";
      s740 <= "0000000000000000000000000000000000";
      s741 <= "0000000000000000000000000000000000";
      s742 <= "0000000000000000000000000000000000";
      s743 <= "0000000000000000000000000000000000";
      s744 <= "0000000000000000000000000000000000";
      s745 <= "0000000000000000000000000000000000";
      s746 <= "0000000000000000000000000000000000";
      s747 <= "0000000000000000000000000000000000";
      s748 <= "0000000000000000000000000000000000";
      s749 <= "0000000000000000000000000000000000";
      s750 <= "0000000000000000000000000000000000";
      s751 <= "0000000000000000000000000000000000";
      s752 <= "0000000000000000000000000000000000";
      s753 <= "0000000000000000000000000000000000";
      s754 <= "0000000000000000000000000000000000";
      s755 <= "0000000000000000000000000000000000";
      s756 <= "0000000000000000000000000000000000";
      s757 <= "0000000000000000000000000000000000";
      s758 <= "0000000000000000000000000000000000";
      s759 <= "0000000000000000000000000000000000";
      s760 <= "0000000000000000000000000000000000";
      s761 <= "0000000000000000000000000000000000";
      s762 <= "0000000000000000000000000000000000";
      s763 <= "0000000000000000000000000000000000";
      s764 <= "0000000000000000000000000000000000";
      s765 <= "0000000000000000000000000000000000";
      s766 <= "0000000000000000000000000000000000";
      s767 <= "0000000000000000000000000000000000";
      s768 <= "0000000000000000000000000000000000";
      s769 <= "0000000000000000000000000000000000";
      s770 <= "0000000000000000000000000000000000";
      s771 <= "0000000000000000000000000000000000";
      s772 <= "0000000000000000000000000000000000";
      s773 <= "0000000000000000000000000000000000";
      s774 <= "0000000000000000000000000000000000";
      s775 <= "0000000000000000000000000000000000";
      s776 <= "0000000000000000000000000000000000";
      s777 <= "0000000000000000000000000000000000";
      s778 <= "0000000000000000000000000000000000";
      s779 <= "0000000000000000000000000000000000";
      s780 <= "0000000000000000000000000000000000";
      s781 <= "0000000000000000000000000000000000";
      s782 <= "0000000000000000000000000000000000";
      s783 <= "0000000000000000000000000000000000";
      s784 <= "0000000000000000000000000000000000";
      s785 <= "0000000000000000000000000000000000";
      s786 <= "0000000000000000000000000000000000";
      s787 <= "0000000000000000000000000000000000";
      s788 <= "0000000000000000000000000000000000";
      s789 <= "0000000000000000000000000000000000";
      s790 <= "0000000000000000000000000000000000";
      s791 <= "0000000000000000000000000000000000";
      s792 <= "0000000000000000000000000000000000";
      s793 <= "0000000000000000000000000000000000";
      s794 <= "0000000000000000000000000000000000";
      s795 <= "0000000000000000000000000000000000";
      s796 <= "0000000000000000000000000000000000";
      s797 <= "0000000000000000000000000000000000";
      s798 <= "0000000000000000000000000000000000";
      s799 <= "0000000000000000000000000000000000";
      s800 <= "0000000000000000000000000000000000";
      s801 <= "0000000000000000000000000000000000";
      s802 <= "0000000000000000000000000000000000";
      s803 <= "0000000000000000000000000000000000";
      s804 <= "0000000000000000000000000000000000";
      s805 <= "0000000000000000000000000000000000";
      s806 <= "0000000000000000000000000000000000";
      s807 <= "0000000000000000000000000000000000";
      s808 <= "0000000000000000000000000000000000";
      s809 <= "0000000000000000000000000000000000";
      s810 <= "0000000000000000000000000000000000";
      s811 <= "0000000000000000000000000000000000";
      s812 <= "0000000000000000000000000000000000";
      s813 <= "0000000000000000000000000000000000";
      s814 <= "0000000000000000000000000000000000";
      s815 <= "0000000000000000000000000000000000";
      s816 <= "0000000000000000000000000000000000";
      s817 <= "0000000000000000000000000000000000";
      s818 <= "0000000000000000000000000000000000";
      s819 <= "0000000000000000000000000000000000";
      s820 <= "0000000000000000000000000000000000";
      s821 <= "0000000000000000000000000000000000";
      s822 <= "0000000000000000000000000000000000";
      s823 <= "0000000000000000000000000000000000";
      s824 <= "0000000000000000000000000000000000";
      s825 <= "0000000000000000000000000000000000";
      s826 <= "0000000000000000000000000000000000";
      s827 <= "0000000000000000000000000000000000";
      s828 <= "0000000000000000000000000000000000";
      s829 <= "0000000000000000000000000000000000";
      s830 <= "0000000000000000000000000000000000";
      s831 <= "0000000000000000000000000000000000";
      s832 <= "0000000000000000000000000000000000";
      s833 <= "0000000000000000000000000000000000";
      s834 <= "0000000000000000000000000000000000";
      s835 <= "0000000000000000000000000000000000";
      s836 <= "0000000000000000000000000000000000";
      s837 <= "0000000000000000000000000000000000";
      s838 <= "0000000000000000000000000000000000";
      s839 <= "0000000000000000000000000000000000";
      s840 <= "0000000000000000000000000000000000";
      s841 <= "0000000000000000000000000000000000";
      s842 <= "0000000000000000000000000000000000";
      s843 <= "0000000000000000000000000000000000";
      s844 <= "0000000000000000000000000000000000";
      s845 <= "0000000000000000000000000000000000";
      s846 <= "0000000000000000000000000000000000";
      s847 <= "0000000000000000000000000000000000";
      s848 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      s558 <= s557;
      s559 <= s558;
      s560 <= s559;
      s561 <= s560;
      s562 <= s561;
      s563 <= s562;
      s564 <= s563;
      s565 <= s564;
      s566 <= s565;
      s567 <= s566;
      s568 <= s567;
      s569 <= s568;
      s570 <= s569;
      s571 <= s570;
      s572 <= s571;
      s573 <= s572;
      s574 <= s573;
      s575 <= s574;
      s576 <= s575;
      s577 <= s576;
      s578 <= s577;
      s579 <= s578;
      s580 <= s579;
      s581 <= s580;
      s582 <= s581;
      s583 <= s582;
      s584 <= s583;
      s585 <= s584;
      s586 <= s585;
      s587 <= s586;
      s588 <= s587;
      s589 <= s588;
      s590 <= s589;
      s591 <= s590;
      s592 <= s591;
      s593 <= s592;
      s594 <= s593;
      s595 <= s594;
      s596 <= s595;
      s597 <= s596;
      s598 <= s597;
      s599 <= s598;
      s600 <= s599;
      s601 <= s600;
      s602 <= s601;
      s603 <= s602;
      s604 <= s603;
      s605 <= s604;
      s606 <= s605;
      s607 <= s606;
      s608 <= s607;
      s609 <= s608;
      s610 <= s609;
      s611 <= s610;
      s612 <= s611;
      s613 <= s612;
      s614 <= s613;
      s615 <= s614;
      s616 <= s615;
      s617 <= s616;
      s618 <= s617;
      s619 <= s618;
      s620 <= s619;
      s621 <= s620;
      s622 <= s621;
      s623 <= s622;
      s624 <= s623;
      s625 <= s624;
      s626 <= s625;
      s627 <= s626;
      s628 <= s627;
      s629 <= s628;
      s630 <= s629;
      s631 <= s630;
      s632 <= s631;
      s633 <= s632;
      s634 <= s633;
      s635 <= s634;
      s636 <= s635;
      s637 <= s636;
      s638 <= s637;
      s639 <= s638;
      s640 <= s639;
      s641 <= s640;
      s642 <= s641;
      s643 <= s642;
      s644 <= s643;
      s645 <= s644;
      s646 <= s645;
      s647 <= s646;
      s648 <= s647;
      s649 <= s648;
      s650 <= s649;
      s651 <= s650;
      s652 <= s651;
      s653 <= s652;
      s654 <= s653;
      s655 <= s654;
      s656 <= s655;
      s657 <= s656;
      s658 <= s657;
      s659 <= s658;
      s660 <= s659;
      s661 <= s660;
      s662 <= s661;
      s663 <= s662;
      s664 <= s663;
      s665 <= s664;
      s666 <= s665;
      s667 <= s666;
      s668 <= s667;
      s669 <= s668;
      s670 <= s669;
      s671 <= s670;
      s672 <= s671;
      s673 <= s672;
      s674 <= s673;
      s675 <= s674;
      s676 <= s675;
      s677 <= s676;
      s678 <= s677;
      s679 <= s678;
      s680 <= s679;
      s681 <= s680;
      s682 <= s681;
      s683 <= s682;
      s684 <= s683;
      s685 <= s684;
      s686 <= s685;
      s687 <= s686;
      s688 <= s687;
      s689 <= s688;
      s690 <= s689;
      s691 <= s690;
      s692 <= s691;
      s693 <= s692;
      s694 <= s693;
      s695 <= s694;
      s696 <= s695;
      s697 <= s696;
      s698 <= s697;
      s699 <= s698;
      s700 <= s699;
      s701 <= s700;
      s702 <= s701;
      s703 <= s702;
      s704 <= s703;
      s705 <= s704;
      s706 <= s705;
      s707 <= s706;
      s708 <= s707;
      s709 <= s708;
      s710 <= s709;
      s711 <= s710;
      s712 <= s711;
      s713 <= s712;
      s714 <= s713;
      s715 <= s714;
      s716 <= s715;
      s717 <= s716;
      s718 <= s717;
      s719 <= s718;
      s720 <= s719;
      s721 <= s720;
      s722 <= s721;
      s723 <= s722;
      s724 <= s723;
      s725 <= s724;
      s726 <= s725;
      s727 <= s726;
      s728 <= s727;
      s729 <= s728;
      s730 <= s729;
      s731 <= s730;
      s732 <= s731;
      s733 <= s732;
      s734 <= s733;
      s735 <= s734;
      s736 <= s735;
      s737 <= s736;
      s738 <= s737;
      s739 <= s738;
      s740 <= s739;
      s741 <= s740;
      s742 <= s741;
      s743 <= s742;
      s744 <= s743;
      s745 <= s744;
      s746 <= s745;
      s747 <= s746;
      s748 <= s747;
      s749 <= s748;
      s750 <= s749;
      s751 <= s750;
      s752 <= s751;
      s753 <= s752;
      s754 <= s753;
      s755 <= s754;
      s756 <= s755;
      s757 <= s756;
      s758 <= s757;
      s759 <= s758;
      s760 <= s759;
      s761 <= s760;
      s762 <= s761;
      s763 <= s762;
      s764 <= s763;
      s765 <= s764;
      s766 <= s765;
      s767 <= s766;
      s768 <= s767;
      s769 <= s768;
      s770 <= s769;
      s771 <= s770;
      s772 <= s771;
      s773 <= s772;
      s774 <= s773;
      s775 <= s774;
      s776 <= s775;
      s777 <= s776;
      s778 <= s777;
      s779 <= s778;
      s780 <= s779;
      s781 <= s780;
      s782 <= s781;
      s783 <= s782;
      s784 <= s783;
      s785 <= s784;
      s786 <= s785;
      s787 <= s786;
      s788 <= s787;
      s789 <= s788;
      s790 <= s789;
      s791 <= s790;
      s792 <= s791;
      s793 <= s792;
      s794 <= s793;
      s795 <= s794;
      s796 <= s795;
      s797 <= s796;
      s798 <= s797;
      s799 <= s798;
      s800 <= s799;
      s801 <= s800;
      s802 <= s801;
      s803 <= s802;
      s804 <= s803;
      s805 <= s804;
      s806 <= s805;
      s807 <= s806;
      s808 <= s807;
      s809 <= s808;
      s810 <= s809;
      s811 <= s810;
      s812 <= s811;
      s813 <= s812;
      s814 <= s813;
      s815 <= s814;
      s816 <= s815;
      s817 <= s816;
      s818 <= s817;
      s819 <= s818;
      s820 <= s819;
      s821 <= s820;
      s822 <= s821;
      s823 <= s822;
      s824 <= s823;
      s825 <= s824;
      s826 <= s825;
      s827 <= s826;
      s828 <= s827;
      s829 <= s828;
      s830 <= s829;
      s831 <= s830;
      s832 <= s831;
      s833 <= s832;
      s834 <= s833;
      s835 <= s834;
      s836 <= s835;
      s837 <= s836;
      s838 <= s837;
      s839 <= s838;
      s840 <= s839;
      s841 <= s840;
      s842 <= s841;
      s843 <= s842;
      s844 <= s843;
      s845 <= s844;
      s846 <= s845;
      s847 <= s846;
      s848 <= s847;
      Y <= s848;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_948_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 948 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_948_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_948_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
signal s558 : std_logic_vector(33 downto 0) := (others => '0');
signal s559 : std_logic_vector(33 downto 0) := (others => '0');
signal s560 : std_logic_vector(33 downto 0) := (others => '0');
signal s561 : std_logic_vector(33 downto 0) := (others => '0');
signal s562 : std_logic_vector(33 downto 0) := (others => '0');
signal s563 : std_logic_vector(33 downto 0) := (others => '0');
signal s564 : std_logic_vector(33 downto 0) := (others => '0');
signal s565 : std_logic_vector(33 downto 0) := (others => '0');
signal s566 : std_logic_vector(33 downto 0) := (others => '0');
signal s567 : std_logic_vector(33 downto 0) := (others => '0');
signal s568 : std_logic_vector(33 downto 0) := (others => '0');
signal s569 : std_logic_vector(33 downto 0) := (others => '0');
signal s570 : std_logic_vector(33 downto 0) := (others => '0');
signal s571 : std_logic_vector(33 downto 0) := (others => '0');
signal s572 : std_logic_vector(33 downto 0) := (others => '0');
signal s573 : std_logic_vector(33 downto 0) := (others => '0');
signal s574 : std_logic_vector(33 downto 0) := (others => '0');
signal s575 : std_logic_vector(33 downto 0) := (others => '0');
signal s576 : std_logic_vector(33 downto 0) := (others => '0');
signal s577 : std_logic_vector(33 downto 0) := (others => '0');
signal s578 : std_logic_vector(33 downto 0) := (others => '0');
signal s579 : std_logic_vector(33 downto 0) := (others => '0');
signal s580 : std_logic_vector(33 downto 0) := (others => '0');
signal s581 : std_logic_vector(33 downto 0) := (others => '0');
signal s582 : std_logic_vector(33 downto 0) := (others => '0');
signal s583 : std_logic_vector(33 downto 0) := (others => '0');
signal s584 : std_logic_vector(33 downto 0) := (others => '0');
signal s585 : std_logic_vector(33 downto 0) := (others => '0');
signal s586 : std_logic_vector(33 downto 0) := (others => '0');
signal s587 : std_logic_vector(33 downto 0) := (others => '0');
signal s588 : std_logic_vector(33 downto 0) := (others => '0');
signal s589 : std_logic_vector(33 downto 0) := (others => '0');
signal s590 : std_logic_vector(33 downto 0) := (others => '0');
signal s591 : std_logic_vector(33 downto 0) := (others => '0');
signal s592 : std_logic_vector(33 downto 0) := (others => '0');
signal s593 : std_logic_vector(33 downto 0) := (others => '0');
signal s594 : std_logic_vector(33 downto 0) := (others => '0');
signal s595 : std_logic_vector(33 downto 0) := (others => '0');
signal s596 : std_logic_vector(33 downto 0) := (others => '0');
signal s597 : std_logic_vector(33 downto 0) := (others => '0');
signal s598 : std_logic_vector(33 downto 0) := (others => '0');
signal s599 : std_logic_vector(33 downto 0) := (others => '0');
signal s600 : std_logic_vector(33 downto 0) := (others => '0');
signal s601 : std_logic_vector(33 downto 0) := (others => '0');
signal s602 : std_logic_vector(33 downto 0) := (others => '0');
signal s603 : std_logic_vector(33 downto 0) := (others => '0');
signal s604 : std_logic_vector(33 downto 0) := (others => '0');
signal s605 : std_logic_vector(33 downto 0) := (others => '0');
signal s606 : std_logic_vector(33 downto 0) := (others => '0');
signal s607 : std_logic_vector(33 downto 0) := (others => '0');
signal s608 : std_logic_vector(33 downto 0) := (others => '0');
signal s609 : std_logic_vector(33 downto 0) := (others => '0');
signal s610 : std_logic_vector(33 downto 0) := (others => '0');
signal s611 : std_logic_vector(33 downto 0) := (others => '0');
signal s612 : std_logic_vector(33 downto 0) := (others => '0');
signal s613 : std_logic_vector(33 downto 0) := (others => '0');
signal s614 : std_logic_vector(33 downto 0) := (others => '0');
signal s615 : std_logic_vector(33 downto 0) := (others => '0');
signal s616 : std_logic_vector(33 downto 0) := (others => '0');
signal s617 : std_logic_vector(33 downto 0) := (others => '0');
signal s618 : std_logic_vector(33 downto 0) := (others => '0');
signal s619 : std_logic_vector(33 downto 0) := (others => '0');
signal s620 : std_logic_vector(33 downto 0) := (others => '0');
signal s621 : std_logic_vector(33 downto 0) := (others => '0');
signal s622 : std_logic_vector(33 downto 0) := (others => '0');
signal s623 : std_logic_vector(33 downto 0) := (others => '0');
signal s624 : std_logic_vector(33 downto 0) := (others => '0');
signal s625 : std_logic_vector(33 downto 0) := (others => '0');
signal s626 : std_logic_vector(33 downto 0) := (others => '0');
signal s627 : std_logic_vector(33 downto 0) := (others => '0');
signal s628 : std_logic_vector(33 downto 0) := (others => '0');
signal s629 : std_logic_vector(33 downto 0) := (others => '0');
signal s630 : std_logic_vector(33 downto 0) := (others => '0');
signal s631 : std_logic_vector(33 downto 0) := (others => '0');
signal s632 : std_logic_vector(33 downto 0) := (others => '0');
signal s633 : std_logic_vector(33 downto 0) := (others => '0');
signal s634 : std_logic_vector(33 downto 0) := (others => '0');
signal s635 : std_logic_vector(33 downto 0) := (others => '0');
signal s636 : std_logic_vector(33 downto 0) := (others => '0');
signal s637 : std_logic_vector(33 downto 0) := (others => '0');
signal s638 : std_logic_vector(33 downto 0) := (others => '0');
signal s639 : std_logic_vector(33 downto 0) := (others => '0');
signal s640 : std_logic_vector(33 downto 0) := (others => '0');
signal s641 : std_logic_vector(33 downto 0) := (others => '0');
signal s642 : std_logic_vector(33 downto 0) := (others => '0');
signal s643 : std_logic_vector(33 downto 0) := (others => '0');
signal s644 : std_logic_vector(33 downto 0) := (others => '0');
signal s645 : std_logic_vector(33 downto 0) := (others => '0');
signal s646 : std_logic_vector(33 downto 0) := (others => '0');
signal s647 : std_logic_vector(33 downto 0) := (others => '0');
signal s648 : std_logic_vector(33 downto 0) := (others => '0');
signal s649 : std_logic_vector(33 downto 0) := (others => '0');
signal s650 : std_logic_vector(33 downto 0) := (others => '0');
signal s651 : std_logic_vector(33 downto 0) := (others => '0');
signal s652 : std_logic_vector(33 downto 0) := (others => '0');
signal s653 : std_logic_vector(33 downto 0) := (others => '0');
signal s654 : std_logic_vector(33 downto 0) := (others => '0');
signal s655 : std_logic_vector(33 downto 0) := (others => '0');
signal s656 : std_logic_vector(33 downto 0) := (others => '0');
signal s657 : std_logic_vector(33 downto 0) := (others => '0');
signal s658 : std_logic_vector(33 downto 0) := (others => '0');
signal s659 : std_logic_vector(33 downto 0) := (others => '0');
signal s660 : std_logic_vector(33 downto 0) := (others => '0');
signal s661 : std_logic_vector(33 downto 0) := (others => '0');
signal s662 : std_logic_vector(33 downto 0) := (others => '0');
signal s663 : std_logic_vector(33 downto 0) := (others => '0');
signal s664 : std_logic_vector(33 downto 0) := (others => '0');
signal s665 : std_logic_vector(33 downto 0) := (others => '0');
signal s666 : std_logic_vector(33 downto 0) := (others => '0');
signal s667 : std_logic_vector(33 downto 0) := (others => '0');
signal s668 : std_logic_vector(33 downto 0) := (others => '0');
signal s669 : std_logic_vector(33 downto 0) := (others => '0');
signal s670 : std_logic_vector(33 downto 0) := (others => '0');
signal s671 : std_logic_vector(33 downto 0) := (others => '0');
signal s672 : std_logic_vector(33 downto 0) := (others => '0');
signal s673 : std_logic_vector(33 downto 0) := (others => '0');
signal s674 : std_logic_vector(33 downto 0) := (others => '0');
signal s675 : std_logic_vector(33 downto 0) := (others => '0');
signal s676 : std_logic_vector(33 downto 0) := (others => '0');
signal s677 : std_logic_vector(33 downto 0) := (others => '0');
signal s678 : std_logic_vector(33 downto 0) := (others => '0');
signal s679 : std_logic_vector(33 downto 0) := (others => '0');
signal s680 : std_logic_vector(33 downto 0) := (others => '0');
signal s681 : std_logic_vector(33 downto 0) := (others => '0');
signal s682 : std_logic_vector(33 downto 0) := (others => '0');
signal s683 : std_logic_vector(33 downto 0) := (others => '0');
signal s684 : std_logic_vector(33 downto 0) := (others => '0');
signal s685 : std_logic_vector(33 downto 0) := (others => '0');
signal s686 : std_logic_vector(33 downto 0) := (others => '0');
signal s687 : std_logic_vector(33 downto 0) := (others => '0');
signal s688 : std_logic_vector(33 downto 0) := (others => '0');
signal s689 : std_logic_vector(33 downto 0) := (others => '0');
signal s690 : std_logic_vector(33 downto 0) := (others => '0');
signal s691 : std_logic_vector(33 downto 0) := (others => '0');
signal s692 : std_logic_vector(33 downto 0) := (others => '0');
signal s693 : std_logic_vector(33 downto 0) := (others => '0');
signal s694 : std_logic_vector(33 downto 0) := (others => '0');
signal s695 : std_logic_vector(33 downto 0) := (others => '0');
signal s696 : std_logic_vector(33 downto 0) := (others => '0');
signal s697 : std_logic_vector(33 downto 0) := (others => '0');
signal s698 : std_logic_vector(33 downto 0) := (others => '0');
signal s699 : std_logic_vector(33 downto 0) := (others => '0');
signal s700 : std_logic_vector(33 downto 0) := (others => '0');
signal s701 : std_logic_vector(33 downto 0) := (others => '0');
signal s702 : std_logic_vector(33 downto 0) := (others => '0');
signal s703 : std_logic_vector(33 downto 0) := (others => '0');
signal s704 : std_logic_vector(33 downto 0) := (others => '0');
signal s705 : std_logic_vector(33 downto 0) := (others => '0');
signal s706 : std_logic_vector(33 downto 0) := (others => '0');
signal s707 : std_logic_vector(33 downto 0) := (others => '0');
signal s708 : std_logic_vector(33 downto 0) := (others => '0');
signal s709 : std_logic_vector(33 downto 0) := (others => '0');
signal s710 : std_logic_vector(33 downto 0) := (others => '0');
signal s711 : std_logic_vector(33 downto 0) := (others => '0');
signal s712 : std_logic_vector(33 downto 0) := (others => '0');
signal s713 : std_logic_vector(33 downto 0) := (others => '0');
signal s714 : std_logic_vector(33 downto 0) := (others => '0');
signal s715 : std_logic_vector(33 downto 0) := (others => '0');
signal s716 : std_logic_vector(33 downto 0) := (others => '0');
signal s717 : std_logic_vector(33 downto 0) := (others => '0');
signal s718 : std_logic_vector(33 downto 0) := (others => '0');
signal s719 : std_logic_vector(33 downto 0) := (others => '0');
signal s720 : std_logic_vector(33 downto 0) := (others => '0');
signal s721 : std_logic_vector(33 downto 0) := (others => '0');
signal s722 : std_logic_vector(33 downto 0) := (others => '0');
signal s723 : std_logic_vector(33 downto 0) := (others => '0');
signal s724 : std_logic_vector(33 downto 0) := (others => '0');
signal s725 : std_logic_vector(33 downto 0) := (others => '0');
signal s726 : std_logic_vector(33 downto 0) := (others => '0');
signal s727 : std_logic_vector(33 downto 0) := (others => '0');
signal s728 : std_logic_vector(33 downto 0) := (others => '0');
signal s729 : std_logic_vector(33 downto 0) := (others => '0');
signal s730 : std_logic_vector(33 downto 0) := (others => '0');
signal s731 : std_logic_vector(33 downto 0) := (others => '0');
signal s732 : std_logic_vector(33 downto 0) := (others => '0');
signal s733 : std_logic_vector(33 downto 0) := (others => '0');
signal s734 : std_logic_vector(33 downto 0) := (others => '0');
signal s735 : std_logic_vector(33 downto 0) := (others => '0');
signal s736 : std_logic_vector(33 downto 0) := (others => '0');
signal s737 : std_logic_vector(33 downto 0) := (others => '0');
signal s738 : std_logic_vector(33 downto 0) := (others => '0');
signal s739 : std_logic_vector(33 downto 0) := (others => '0');
signal s740 : std_logic_vector(33 downto 0) := (others => '0');
signal s741 : std_logic_vector(33 downto 0) := (others => '0');
signal s742 : std_logic_vector(33 downto 0) := (others => '0');
signal s743 : std_logic_vector(33 downto 0) := (others => '0');
signal s744 : std_logic_vector(33 downto 0) := (others => '0');
signal s745 : std_logic_vector(33 downto 0) := (others => '0');
signal s746 : std_logic_vector(33 downto 0) := (others => '0');
signal s747 : std_logic_vector(33 downto 0) := (others => '0');
signal s748 : std_logic_vector(33 downto 0) := (others => '0');
signal s749 : std_logic_vector(33 downto 0) := (others => '0');
signal s750 : std_logic_vector(33 downto 0) := (others => '0');
signal s751 : std_logic_vector(33 downto 0) := (others => '0');
signal s752 : std_logic_vector(33 downto 0) := (others => '0');
signal s753 : std_logic_vector(33 downto 0) := (others => '0');
signal s754 : std_logic_vector(33 downto 0) := (others => '0');
signal s755 : std_logic_vector(33 downto 0) := (others => '0');
signal s756 : std_logic_vector(33 downto 0) := (others => '0');
signal s757 : std_logic_vector(33 downto 0) := (others => '0');
signal s758 : std_logic_vector(33 downto 0) := (others => '0');
signal s759 : std_logic_vector(33 downto 0) := (others => '0');
signal s760 : std_logic_vector(33 downto 0) := (others => '0');
signal s761 : std_logic_vector(33 downto 0) := (others => '0');
signal s762 : std_logic_vector(33 downto 0) := (others => '0');
signal s763 : std_logic_vector(33 downto 0) := (others => '0');
signal s764 : std_logic_vector(33 downto 0) := (others => '0');
signal s765 : std_logic_vector(33 downto 0) := (others => '0');
signal s766 : std_logic_vector(33 downto 0) := (others => '0');
signal s767 : std_logic_vector(33 downto 0) := (others => '0');
signal s768 : std_logic_vector(33 downto 0) := (others => '0');
signal s769 : std_logic_vector(33 downto 0) := (others => '0');
signal s770 : std_logic_vector(33 downto 0) := (others => '0');
signal s771 : std_logic_vector(33 downto 0) := (others => '0');
signal s772 : std_logic_vector(33 downto 0) := (others => '0');
signal s773 : std_logic_vector(33 downto 0) := (others => '0');
signal s774 : std_logic_vector(33 downto 0) := (others => '0');
signal s775 : std_logic_vector(33 downto 0) := (others => '0');
signal s776 : std_logic_vector(33 downto 0) := (others => '0');
signal s777 : std_logic_vector(33 downto 0) := (others => '0');
signal s778 : std_logic_vector(33 downto 0) := (others => '0');
signal s779 : std_logic_vector(33 downto 0) := (others => '0');
signal s780 : std_logic_vector(33 downto 0) := (others => '0');
signal s781 : std_logic_vector(33 downto 0) := (others => '0');
signal s782 : std_logic_vector(33 downto 0) := (others => '0');
signal s783 : std_logic_vector(33 downto 0) := (others => '0');
signal s784 : std_logic_vector(33 downto 0) := (others => '0');
signal s785 : std_logic_vector(33 downto 0) := (others => '0');
signal s786 : std_logic_vector(33 downto 0) := (others => '0');
signal s787 : std_logic_vector(33 downto 0) := (others => '0');
signal s788 : std_logic_vector(33 downto 0) := (others => '0');
signal s789 : std_logic_vector(33 downto 0) := (others => '0');
signal s790 : std_logic_vector(33 downto 0) := (others => '0');
signal s791 : std_logic_vector(33 downto 0) := (others => '0');
signal s792 : std_logic_vector(33 downto 0) := (others => '0');
signal s793 : std_logic_vector(33 downto 0) := (others => '0');
signal s794 : std_logic_vector(33 downto 0) := (others => '0');
signal s795 : std_logic_vector(33 downto 0) := (others => '0');
signal s796 : std_logic_vector(33 downto 0) := (others => '0');
signal s797 : std_logic_vector(33 downto 0) := (others => '0');
signal s798 : std_logic_vector(33 downto 0) := (others => '0');
signal s799 : std_logic_vector(33 downto 0) := (others => '0');
signal s800 : std_logic_vector(33 downto 0) := (others => '0');
signal s801 : std_logic_vector(33 downto 0) := (others => '0');
signal s802 : std_logic_vector(33 downto 0) := (others => '0');
signal s803 : std_logic_vector(33 downto 0) := (others => '0');
signal s804 : std_logic_vector(33 downto 0) := (others => '0');
signal s805 : std_logic_vector(33 downto 0) := (others => '0');
signal s806 : std_logic_vector(33 downto 0) := (others => '0');
signal s807 : std_logic_vector(33 downto 0) := (others => '0');
signal s808 : std_logic_vector(33 downto 0) := (others => '0');
signal s809 : std_logic_vector(33 downto 0) := (others => '0');
signal s810 : std_logic_vector(33 downto 0) := (others => '0');
signal s811 : std_logic_vector(33 downto 0) := (others => '0');
signal s812 : std_logic_vector(33 downto 0) := (others => '0');
signal s813 : std_logic_vector(33 downto 0) := (others => '0');
signal s814 : std_logic_vector(33 downto 0) := (others => '0');
signal s815 : std_logic_vector(33 downto 0) := (others => '0');
signal s816 : std_logic_vector(33 downto 0) := (others => '0');
signal s817 : std_logic_vector(33 downto 0) := (others => '0');
signal s818 : std_logic_vector(33 downto 0) := (others => '0');
signal s819 : std_logic_vector(33 downto 0) := (others => '0');
signal s820 : std_logic_vector(33 downto 0) := (others => '0');
signal s821 : std_logic_vector(33 downto 0) := (others => '0');
signal s822 : std_logic_vector(33 downto 0) := (others => '0');
signal s823 : std_logic_vector(33 downto 0) := (others => '0');
signal s824 : std_logic_vector(33 downto 0) := (others => '0');
signal s825 : std_logic_vector(33 downto 0) := (others => '0');
signal s826 : std_logic_vector(33 downto 0) := (others => '0');
signal s827 : std_logic_vector(33 downto 0) := (others => '0');
signal s828 : std_logic_vector(33 downto 0) := (others => '0');
signal s829 : std_logic_vector(33 downto 0) := (others => '0');
signal s830 : std_logic_vector(33 downto 0) := (others => '0');
signal s831 : std_logic_vector(33 downto 0) := (others => '0');
signal s832 : std_logic_vector(33 downto 0) := (others => '0');
signal s833 : std_logic_vector(33 downto 0) := (others => '0');
signal s834 : std_logic_vector(33 downto 0) := (others => '0');
signal s835 : std_logic_vector(33 downto 0) := (others => '0');
signal s836 : std_logic_vector(33 downto 0) := (others => '0');
signal s837 : std_logic_vector(33 downto 0) := (others => '0');
signal s838 : std_logic_vector(33 downto 0) := (others => '0');
signal s839 : std_logic_vector(33 downto 0) := (others => '0');
signal s840 : std_logic_vector(33 downto 0) := (others => '0');
signal s841 : std_logic_vector(33 downto 0) := (others => '0');
signal s842 : std_logic_vector(33 downto 0) := (others => '0');
signal s843 : std_logic_vector(33 downto 0) := (others => '0');
signal s844 : std_logic_vector(33 downto 0) := (others => '0');
signal s845 : std_logic_vector(33 downto 0) := (others => '0');
signal s846 : std_logic_vector(33 downto 0) := (others => '0');
signal s847 : std_logic_vector(33 downto 0) := (others => '0');
signal s848 : std_logic_vector(33 downto 0) := (others => '0');
signal s849 : std_logic_vector(33 downto 0) := (others => '0');
signal s850 : std_logic_vector(33 downto 0) := (others => '0');
signal s851 : std_logic_vector(33 downto 0) := (others => '0');
signal s852 : std_logic_vector(33 downto 0) := (others => '0');
signal s853 : std_logic_vector(33 downto 0) := (others => '0');
signal s854 : std_logic_vector(33 downto 0) := (others => '0');
signal s855 : std_logic_vector(33 downto 0) := (others => '0');
signal s856 : std_logic_vector(33 downto 0) := (others => '0');
signal s857 : std_logic_vector(33 downto 0) := (others => '0');
signal s858 : std_logic_vector(33 downto 0) := (others => '0');
signal s859 : std_logic_vector(33 downto 0) := (others => '0');
signal s860 : std_logic_vector(33 downto 0) := (others => '0');
signal s861 : std_logic_vector(33 downto 0) := (others => '0');
signal s862 : std_logic_vector(33 downto 0) := (others => '0');
signal s863 : std_logic_vector(33 downto 0) := (others => '0');
signal s864 : std_logic_vector(33 downto 0) := (others => '0');
signal s865 : std_logic_vector(33 downto 0) := (others => '0');
signal s866 : std_logic_vector(33 downto 0) := (others => '0');
signal s867 : std_logic_vector(33 downto 0) := (others => '0');
signal s868 : std_logic_vector(33 downto 0) := (others => '0');
signal s869 : std_logic_vector(33 downto 0) := (others => '0');
signal s870 : std_logic_vector(33 downto 0) := (others => '0');
signal s871 : std_logic_vector(33 downto 0) := (others => '0');
signal s872 : std_logic_vector(33 downto 0) := (others => '0');
signal s873 : std_logic_vector(33 downto 0) := (others => '0');
signal s874 : std_logic_vector(33 downto 0) := (others => '0');
signal s875 : std_logic_vector(33 downto 0) := (others => '0');
signal s876 : std_logic_vector(33 downto 0) := (others => '0');
signal s877 : std_logic_vector(33 downto 0) := (others => '0');
signal s878 : std_logic_vector(33 downto 0) := (others => '0');
signal s879 : std_logic_vector(33 downto 0) := (others => '0');
signal s880 : std_logic_vector(33 downto 0) := (others => '0');
signal s881 : std_logic_vector(33 downto 0) := (others => '0');
signal s882 : std_logic_vector(33 downto 0) := (others => '0');
signal s883 : std_logic_vector(33 downto 0) := (others => '0');
signal s884 : std_logic_vector(33 downto 0) := (others => '0');
signal s885 : std_logic_vector(33 downto 0) := (others => '0');
signal s886 : std_logic_vector(33 downto 0) := (others => '0');
signal s887 : std_logic_vector(33 downto 0) := (others => '0');
signal s888 : std_logic_vector(33 downto 0) := (others => '0');
signal s889 : std_logic_vector(33 downto 0) := (others => '0');
signal s890 : std_logic_vector(33 downto 0) := (others => '0');
signal s891 : std_logic_vector(33 downto 0) := (others => '0');
signal s892 : std_logic_vector(33 downto 0) := (others => '0');
signal s893 : std_logic_vector(33 downto 0) := (others => '0');
signal s894 : std_logic_vector(33 downto 0) := (others => '0');
signal s895 : std_logic_vector(33 downto 0) := (others => '0');
signal s896 : std_logic_vector(33 downto 0) := (others => '0');
signal s897 : std_logic_vector(33 downto 0) := (others => '0');
signal s898 : std_logic_vector(33 downto 0) := (others => '0');
signal s899 : std_logic_vector(33 downto 0) := (others => '0');
signal s900 : std_logic_vector(33 downto 0) := (others => '0');
signal s901 : std_logic_vector(33 downto 0) := (others => '0');
signal s902 : std_logic_vector(33 downto 0) := (others => '0');
signal s903 : std_logic_vector(33 downto 0) := (others => '0');
signal s904 : std_logic_vector(33 downto 0) := (others => '0');
signal s905 : std_logic_vector(33 downto 0) := (others => '0');
signal s906 : std_logic_vector(33 downto 0) := (others => '0');
signal s907 : std_logic_vector(33 downto 0) := (others => '0');
signal s908 : std_logic_vector(33 downto 0) := (others => '0');
signal s909 : std_logic_vector(33 downto 0) := (others => '0');
signal s910 : std_logic_vector(33 downto 0) := (others => '0');
signal s911 : std_logic_vector(33 downto 0) := (others => '0');
signal s912 : std_logic_vector(33 downto 0) := (others => '0');
signal s913 : std_logic_vector(33 downto 0) := (others => '0');
signal s914 : std_logic_vector(33 downto 0) := (others => '0');
signal s915 : std_logic_vector(33 downto 0) := (others => '0');
signal s916 : std_logic_vector(33 downto 0) := (others => '0');
signal s917 : std_logic_vector(33 downto 0) := (others => '0');
signal s918 : std_logic_vector(33 downto 0) := (others => '0');
signal s919 : std_logic_vector(33 downto 0) := (others => '0');
signal s920 : std_logic_vector(33 downto 0) := (others => '0');
signal s921 : std_logic_vector(33 downto 0) := (others => '0');
signal s922 : std_logic_vector(33 downto 0) := (others => '0');
signal s923 : std_logic_vector(33 downto 0) := (others => '0');
signal s924 : std_logic_vector(33 downto 0) := (others => '0');
signal s925 : std_logic_vector(33 downto 0) := (others => '0');
signal s926 : std_logic_vector(33 downto 0) := (others => '0');
signal s927 : std_logic_vector(33 downto 0) := (others => '0');
signal s928 : std_logic_vector(33 downto 0) := (others => '0');
signal s929 : std_logic_vector(33 downto 0) := (others => '0');
signal s930 : std_logic_vector(33 downto 0) := (others => '0');
signal s931 : std_logic_vector(33 downto 0) := (others => '0');
signal s932 : std_logic_vector(33 downto 0) := (others => '0');
signal s933 : std_logic_vector(33 downto 0) := (others => '0');
signal s934 : std_logic_vector(33 downto 0) := (others => '0');
signal s935 : std_logic_vector(33 downto 0) := (others => '0');
signal s936 : std_logic_vector(33 downto 0) := (others => '0');
signal s937 : std_logic_vector(33 downto 0) := (others => '0');
signal s938 : std_logic_vector(33 downto 0) := (others => '0');
signal s939 : std_logic_vector(33 downto 0) := (others => '0');
signal s940 : std_logic_vector(33 downto 0) := (others => '0');
signal s941 : std_logic_vector(33 downto 0) := (others => '0');
signal s942 : std_logic_vector(33 downto 0) := (others => '0');
signal s943 : std_logic_vector(33 downto 0) := (others => '0');
signal s944 : std_logic_vector(33 downto 0) := (others => '0');
signal s945 : std_logic_vector(33 downto 0) := (others => '0');
signal s946 : std_logic_vector(33 downto 0) := (others => '0');
signal s947 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
      s558 <= "0000000000000000000000000000000000";
      s559 <= "0000000000000000000000000000000000";
      s560 <= "0000000000000000000000000000000000";
      s561 <= "0000000000000000000000000000000000";
      s562 <= "0000000000000000000000000000000000";
      s563 <= "0000000000000000000000000000000000";
      s564 <= "0000000000000000000000000000000000";
      s565 <= "0000000000000000000000000000000000";
      s566 <= "0000000000000000000000000000000000";
      s567 <= "0000000000000000000000000000000000";
      s568 <= "0000000000000000000000000000000000";
      s569 <= "0000000000000000000000000000000000";
      s570 <= "0000000000000000000000000000000000";
      s571 <= "0000000000000000000000000000000000";
      s572 <= "0000000000000000000000000000000000";
      s573 <= "0000000000000000000000000000000000";
      s574 <= "0000000000000000000000000000000000";
      s575 <= "0000000000000000000000000000000000";
      s576 <= "0000000000000000000000000000000000";
      s577 <= "0000000000000000000000000000000000";
      s578 <= "0000000000000000000000000000000000";
      s579 <= "0000000000000000000000000000000000";
      s580 <= "0000000000000000000000000000000000";
      s581 <= "0000000000000000000000000000000000";
      s582 <= "0000000000000000000000000000000000";
      s583 <= "0000000000000000000000000000000000";
      s584 <= "0000000000000000000000000000000000";
      s585 <= "0000000000000000000000000000000000";
      s586 <= "0000000000000000000000000000000000";
      s587 <= "0000000000000000000000000000000000";
      s588 <= "0000000000000000000000000000000000";
      s589 <= "0000000000000000000000000000000000";
      s590 <= "0000000000000000000000000000000000";
      s591 <= "0000000000000000000000000000000000";
      s592 <= "0000000000000000000000000000000000";
      s593 <= "0000000000000000000000000000000000";
      s594 <= "0000000000000000000000000000000000";
      s595 <= "0000000000000000000000000000000000";
      s596 <= "0000000000000000000000000000000000";
      s597 <= "0000000000000000000000000000000000";
      s598 <= "0000000000000000000000000000000000";
      s599 <= "0000000000000000000000000000000000";
      s600 <= "0000000000000000000000000000000000";
      s601 <= "0000000000000000000000000000000000";
      s602 <= "0000000000000000000000000000000000";
      s603 <= "0000000000000000000000000000000000";
      s604 <= "0000000000000000000000000000000000";
      s605 <= "0000000000000000000000000000000000";
      s606 <= "0000000000000000000000000000000000";
      s607 <= "0000000000000000000000000000000000";
      s608 <= "0000000000000000000000000000000000";
      s609 <= "0000000000000000000000000000000000";
      s610 <= "0000000000000000000000000000000000";
      s611 <= "0000000000000000000000000000000000";
      s612 <= "0000000000000000000000000000000000";
      s613 <= "0000000000000000000000000000000000";
      s614 <= "0000000000000000000000000000000000";
      s615 <= "0000000000000000000000000000000000";
      s616 <= "0000000000000000000000000000000000";
      s617 <= "0000000000000000000000000000000000";
      s618 <= "0000000000000000000000000000000000";
      s619 <= "0000000000000000000000000000000000";
      s620 <= "0000000000000000000000000000000000";
      s621 <= "0000000000000000000000000000000000";
      s622 <= "0000000000000000000000000000000000";
      s623 <= "0000000000000000000000000000000000";
      s624 <= "0000000000000000000000000000000000";
      s625 <= "0000000000000000000000000000000000";
      s626 <= "0000000000000000000000000000000000";
      s627 <= "0000000000000000000000000000000000";
      s628 <= "0000000000000000000000000000000000";
      s629 <= "0000000000000000000000000000000000";
      s630 <= "0000000000000000000000000000000000";
      s631 <= "0000000000000000000000000000000000";
      s632 <= "0000000000000000000000000000000000";
      s633 <= "0000000000000000000000000000000000";
      s634 <= "0000000000000000000000000000000000";
      s635 <= "0000000000000000000000000000000000";
      s636 <= "0000000000000000000000000000000000";
      s637 <= "0000000000000000000000000000000000";
      s638 <= "0000000000000000000000000000000000";
      s639 <= "0000000000000000000000000000000000";
      s640 <= "0000000000000000000000000000000000";
      s641 <= "0000000000000000000000000000000000";
      s642 <= "0000000000000000000000000000000000";
      s643 <= "0000000000000000000000000000000000";
      s644 <= "0000000000000000000000000000000000";
      s645 <= "0000000000000000000000000000000000";
      s646 <= "0000000000000000000000000000000000";
      s647 <= "0000000000000000000000000000000000";
      s648 <= "0000000000000000000000000000000000";
      s649 <= "0000000000000000000000000000000000";
      s650 <= "0000000000000000000000000000000000";
      s651 <= "0000000000000000000000000000000000";
      s652 <= "0000000000000000000000000000000000";
      s653 <= "0000000000000000000000000000000000";
      s654 <= "0000000000000000000000000000000000";
      s655 <= "0000000000000000000000000000000000";
      s656 <= "0000000000000000000000000000000000";
      s657 <= "0000000000000000000000000000000000";
      s658 <= "0000000000000000000000000000000000";
      s659 <= "0000000000000000000000000000000000";
      s660 <= "0000000000000000000000000000000000";
      s661 <= "0000000000000000000000000000000000";
      s662 <= "0000000000000000000000000000000000";
      s663 <= "0000000000000000000000000000000000";
      s664 <= "0000000000000000000000000000000000";
      s665 <= "0000000000000000000000000000000000";
      s666 <= "0000000000000000000000000000000000";
      s667 <= "0000000000000000000000000000000000";
      s668 <= "0000000000000000000000000000000000";
      s669 <= "0000000000000000000000000000000000";
      s670 <= "0000000000000000000000000000000000";
      s671 <= "0000000000000000000000000000000000";
      s672 <= "0000000000000000000000000000000000";
      s673 <= "0000000000000000000000000000000000";
      s674 <= "0000000000000000000000000000000000";
      s675 <= "0000000000000000000000000000000000";
      s676 <= "0000000000000000000000000000000000";
      s677 <= "0000000000000000000000000000000000";
      s678 <= "0000000000000000000000000000000000";
      s679 <= "0000000000000000000000000000000000";
      s680 <= "0000000000000000000000000000000000";
      s681 <= "0000000000000000000000000000000000";
      s682 <= "0000000000000000000000000000000000";
      s683 <= "0000000000000000000000000000000000";
      s684 <= "0000000000000000000000000000000000";
      s685 <= "0000000000000000000000000000000000";
      s686 <= "0000000000000000000000000000000000";
      s687 <= "0000000000000000000000000000000000";
      s688 <= "0000000000000000000000000000000000";
      s689 <= "0000000000000000000000000000000000";
      s690 <= "0000000000000000000000000000000000";
      s691 <= "0000000000000000000000000000000000";
      s692 <= "0000000000000000000000000000000000";
      s693 <= "0000000000000000000000000000000000";
      s694 <= "0000000000000000000000000000000000";
      s695 <= "0000000000000000000000000000000000";
      s696 <= "0000000000000000000000000000000000";
      s697 <= "0000000000000000000000000000000000";
      s698 <= "0000000000000000000000000000000000";
      s699 <= "0000000000000000000000000000000000";
      s700 <= "0000000000000000000000000000000000";
      s701 <= "0000000000000000000000000000000000";
      s702 <= "0000000000000000000000000000000000";
      s703 <= "0000000000000000000000000000000000";
      s704 <= "0000000000000000000000000000000000";
      s705 <= "0000000000000000000000000000000000";
      s706 <= "0000000000000000000000000000000000";
      s707 <= "0000000000000000000000000000000000";
      s708 <= "0000000000000000000000000000000000";
      s709 <= "0000000000000000000000000000000000";
      s710 <= "0000000000000000000000000000000000";
      s711 <= "0000000000000000000000000000000000";
      s712 <= "0000000000000000000000000000000000";
      s713 <= "0000000000000000000000000000000000";
      s714 <= "0000000000000000000000000000000000";
      s715 <= "0000000000000000000000000000000000";
      s716 <= "0000000000000000000000000000000000";
      s717 <= "0000000000000000000000000000000000";
      s718 <= "0000000000000000000000000000000000";
      s719 <= "0000000000000000000000000000000000";
      s720 <= "0000000000000000000000000000000000";
      s721 <= "0000000000000000000000000000000000";
      s722 <= "0000000000000000000000000000000000";
      s723 <= "0000000000000000000000000000000000";
      s724 <= "0000000000000000000000000000000000";
      s725 <= "0000000000000000000000000000000000";
      s726 <= "0000000000000000000000000000000000";
      s727 <= "0000000000000000000000000000000000";
      s728 <= "0000000000000000000000000000000000";
      s729 <= "0000000000000000000000000000000000";
      s730 <= "0000000000000000000000000000000000";
      s731 <= "0000000000000000000000000000000000";
      s732 <= "0000000000000000000000000000000000";
      s733 <= "0000000000000000000000000000000000";
      s734 <= "0000000000000000000000000000000000";
      s735 <= "0000000000000000000000000000000000";
      s736 <= "0000000000000000000000000000000000";
      s737 <= "0000000000000000000000000000000000";
      s738 <= "0000000000000000000000000000000000";
      s739 <= "0000000000000000000000000000000000";
      s740 <= "0000000000000000000000000000000000";
      s741 <= "0000000000000000000000000000000000";
      s742 <= "0000000000000000000000000000000000";
      s743 <= "0000000000000000000000000000000000";
      s744 <= "0000000000000000000000000000000000";
      s745 <= "0000000000000000000000000000000000";
      s746 <= "0000000000000000000000000000000000";
      s747 <= "0000000000000000000000000000000000";
      s748 <= "0000000000000000000000000000000000";
      s749 <= "0000000000000000000000000000000000";
      s750 <= "0000000000000000000000000000000000";
      s751 <= "0000000000000000000000000000000000";
      s752 <= "0000000000000000000000000000000000";
      s753 <= "0000000000000000000000000000000000";
      s754 <= "0000000000000000000000000000000000";
      s755 <= "0000000000000000000000000000000000";
      s756 <= "0000000000000000000000000000000000";
      s757 <= "0000000000000000000000000000000000";
      s758 <= "0000000000000000000000000000000000";
      s759 <= "0000000000000000000000000000000000";
      s760 <= "0000000000000000000000000000000000";
      s761 <= "0000000000000000000000000000000000";
      s762 <= "0000000000000000000000000000000000";
      s763 <= "0000000000000000000000000000000000";
      s764 <= "0000000000000000000000000000000000";
      s765 <= "0000000000000000000000000000000000";
      s766 <= "0000000000000000000000000000000000";
      s767 <= "0000000000000000000000000000000000";
      s768 <= "0000000000000000000000000000000000";
      s769 <= "0000000000000000000000000000000000";
      s770 <= "0000000000000000000000000000000000";
      s771 <= "0000000000000000000000000000000000";
      s772 <= "0000000000000000000000000000000000";
      s773 <= "0000000000000000000000000000000000";
      s774 <= "0000000000000000000000000000000000";
      s775 <= "0000000000000000000000000000000000";
      s776 <= "0000000000000000000000000000000000";
      s777 <= "0000000000000000000000000000000000";
      s778 <= "0000000000000000000000000000000000";
      s779 <= "0000000000000000000000000000000000";
      s780 <= "0000000000000000000000000000000000";
      s781 <= "0000000000000000000000000000000000";
      s782 <= "0000000000000000000000000000000000";
      s783 <= "0000000000000000000000000000000000";
      s784 <= "0000000000000000000000000000000000";
      s785 <= "0000000000000000000000000000000000";
      s786 <= "0000000000000000000000000000000000";
      s787 <= "0000000000000000000000000000000000";
      s788 <= "0000000000000000000000000000000000";
      s789 <= "0000000000000000000000000000000000";
      s790 <= "0000000000000000000000000000000000";
      s791 <= "0000000000000000000000000000000000";
      s792 <= "0000000000000000000000000000000000";
      s793 <= "0000000000000000000000000000000000";
      s794 <= "0000000000000000000000000000000000";
      s795 <= "0000000000000000000000000000000000";
      s796 <= "0000000000000000000000000000000000";
      s797 <= "0000000000000000000000000000000000";
      s798 <= "0000000000000000000000000000000000";
      s799 <= "0000000000000000000000000000000000";
      s800 <= "0000000000000000000000000000000000";
      s801 <= "0000000000000000000000000000000000";
      s802 <= "0000000000000000000000000000000000";
      s803 <= "0000000000000000000000000000000000";
      s804 <= "0000000000000000000000000000000000";
      s805 <= "0000000000000000000000000000000000";
      s806 <= "0000000000000000000000000000000000";
      s807 <= "0000000000000000000000000000000000";
      s808 <= "0000000000000000000000000000000000";
      s809 <= "0000000000000000000000000000000000";
      s810 <= "0000000000000000000000000000000000";
      s811 <= "0000000000000000000000000000000000";
      s812 <= "0000000000000000000000000000000000";
      s813 <= "0000000000000000000000000000000000";
      s814 <= "0000000000000000000000000000000000";
      s815 <= "0000000000000000000000000000000000";
      s816 <= "0000000000000000000000000000000000";
      s817 <= "0000000000000000000000000000000000";
      s818 <= "0000000000000000000000000000000000";
      s819 <= "0000000000000000000000000000000000";
      s820 <= "0000000000000000000000000000000000";
      s821 <= "0000000000000000000000000000000000";
      s822 <= "0000000000000000000000000000000000";
      s823 <= "0000000000000000000000000000000000";
      s824 <= "0000000000000000000000000000000000";
      s825 <= "0000000000000000000000000000000000";
      s826 <= "0000000000000000000000000000000000";
      s827 <= "0000000000000000000000000000000000";
      s828 <= "0000000000000000000000000000000000";
      s829 <= "0000000000000000000000000000000000";
      s830 <= "0000000000000000000000000000000000";
      s831 <= "0000000000000000000000000000000000";
      s832 <= "0000000000000000000000000000000000";
      s833 <= "0000000000000000000000000000000000";
      s834 <= "0000000000000000000000000000000000";
      s835 <= "0000000000000000000000000000000000";
      s836 <= "0000000000000000000000000000000000";
      s837 <= "0000000000000000000000000000000000";
      s838 <= "0000000000000000000000000000000000";
      s839 <= "0000000000000000000000000000000000";
      s840 <= "0000000000000000000000000000000000";
      s841 <= "0000000000000000000000000000000000";
      s842 <= "0000000000000000000000000000000000";
      s843 <= "0000000000000000000000000000000000";
      s844 <= "0000000000000000000000000000000000";
      s845 <= "0000000000000000000000000000000000";
      s846 <= "0000000000000000000000000000000000";
      s847 <= "0000000000000000000000000000000000";
      s848 <= "0000000000000000000000000000000000";
      s849 <= "0000000000000000000000000000000000";
      s850 <= "0000000000000000000000000000000000";
      s851 <= "0000000000000000000000000000000000";
      s852 <= "0000000000000000000000000000000000";
      s853 <= "0000000000000000000000000000000000";
      s854 <= "0000000000000000000000000000000000";
      s855 <= "0000000000000000000000000000000000";
      s856 <= "0000000000000000000000000000000000";
      s857 <= "0000000000000000000000000000000000";
      s858 <= "0000000000000000000000000000000000";
      s859 <= "0000000000000000000000000000000000";
      s860 <= "0000000000000000000000000000000000";
      s861 <= "0000000000000000000000000000000000";
      s862 <= "0000000000000000000000000000000000";
      s863 <= "0000000000000000000000000000000000";
      s864 <= "0000000000000000000000000000000000";
      s865 <= "0000000000000000000000000000000000";
      s866 <= "0000000000000000000000000000000000";
      s867 <= "0000000000000000000000000000000000";
      s868 <= "0000000000000000000000000000000000";
      s869 <= "0000000000000000000000000000000000";
      s870 <= "0000000000000000000000000000000000";
      s871 <= "0000000000000000000000000000000000";
      s872 <= "0000000000000000000000000000000000";
      s873 <= "0000000000000000000000000000000000";
      s874 <= "0000000000000000000000000000000000";
      s875 <= "0000000000000000000000000000000000";
      s876 <= "0000000000000000000000000000000000";
      s877 <= "0000000000000000000000000000000000";
      s878 <= "0000000000000000000000000000000000";
      s879 <= "0000000000000000000000000000000000";
      s880 <= "0000000000000000000000000000000000";
      s881 <= "0000000000000000000000000000000000";
      s882 <= "0000000000000000000000000000000000";
      s883 <= "0000000000000000000000000000000000";
      s884 <= "0000000000000000000000000000000000";
      s885 <= "0000000000000000000000000000000000";
      s886 <= "0000000000000000000000000000000000";
      s887 <= "0000000000000000000000000000000000";
      s888 <= "0000000000000000000000000000000000";
      s889 <= "0000000000000000000000000000000000";
      s890 <= "0000000000000000000000000000000000";
      s891 <= "0000000000000000000000000000000000";
      s892 <= "0000000000000000000000000000000000";
      s893 <= "0000000000000000000000000000000000";
      s894 <= "0000000000000000000000000000000000";
      s895 <= "0000000000000000000000000000000000";
      s896 <= "0000000000000000000000000000000000";
      s897 <= "0000000000000000000000000000000000";
      s898 <= "0000000000000000000000000000000000";
      s899 <= "0000000000000000000000000000000000";
      s900 <= "0000000000000000000000000000000000";
      s901 <= "0000000000000000000000000000000000";
      s902 <= "0000000000000000000000000000000000";
      s903 <= "0000000000000000000000000000000000";
      s904 <= "0000000000000000000000000000000000";
      s905 <= "0000000000000000000000000000000000";
      s906 <= "0000000000000000000000000000000000";
      s907 <= "0000000000000000000000000000000000";
      s908 <= "0000000000000000000000000000000000";
      s909 <= "0000000000000000000000000000000000";
      s910 <= "0000000000000000000000000000000000";
      s911 <= "0000000000000000000000000000000000";
      s912 <= "0000000000000000000000000000000000";
      s913 <= "0000000000000000000000000000000000";
      s914 <= "0000000000000000000000000000000000";
      s915 <= "0000000000000000000000000000000000";
      s916 <= "0000000000000000000000000000000000";
      s917 <= "0000000000000000000000000000000000";
      s918 <= "0000000000000000000000000000000000";
      s919 <= "0000000000000000000000000000000000";
      s920 <= "0000000000000000000000000000000000";
      s921 <= "0000000000000000000000000000000000";
      s922 <= "0000000000000000000000000000000000";
      s923 <= "0000000000000000000000000000000000";
      s924 <= "0000000000000000000000000000000000";
      s925 <= "0000000000000000000000000000000000";
      s926 <= "0000000000000000000000000000000000";
      s927 <= "0000000000000000000000000000000000";
      s928 <= "0000000000000000000000000000000000";
      s929 <= "0000000000000000000000000000000000";
      s930 <= "0000000000000000000000000000000000";
      s931 <= "0000000000000000000000000000000000";
      s932 <= "0000000000000000000000000000000000";
      s933 <= "0000000000000000000000000000000000";
      s934 <= "0000000000000000000000000000000000";
      s935 <= "0000000000000000000000000000000000";
      s936 <= "0000000000000000000000000000000000";
      s937 <= "0000000000000000000000000000000000";
      s938 <= "0000000000000000000000000000000000";
      s939 <= "0000000000000000000000000000000000";
      s940 <= "0000000000000000000000000000000000";
      s941 <= "0000000000000000000000000000000000";
      s942 <= "0000000000000000000000000000000000";
      s943 <= "0000000000000000000000000000000000";
      s944 <= "0000000000000000000000000000000000";
      s945 <= "0000000000000000000000000000000000";
      s946 <= "0000000000000000000000000000000000";
      s947 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      s558 <= s557;
      s559 <= s558;
      s560 <= s559;
      s561 <= s560;
      s562 <= s561;
      s563 <= s562;
      s564 <= s563;
      s565 <= s564;
      s566 <= s565;
      s567 <= s566;
      s568 <= s567;
      s569 <= s568;
      s570 <= s569;
      s571 <= s570;
      s572 <= s571;
      s573 <= s572;
      s574 <= s573;
      s575 <= s574;
      s576 <= s575;
      s577 <= s576;
      s578 <= s577;
      s579 <= s578;
      s580 <= s579;
      s581 <= s580;
      s582 <= s581;
      s583 <= s582;
      s584 <= s583;
      s585 <= s584;
      s586 <= s585;
      s587 <= s586;
      s588 <= s587;
      s589 <= s588;
      s590 <= s589;
      s591 <= s590;
      s592 <= s591;
      s593 <= s592;
      s594 <= s593;
      s595 <= s594;
      s596 <= s595;
      s597 <= s596;
      s598 <= s597;
      s599 <= s598;
      s600 <= s599;
      s601 <= s600;
      s602 <= s601;
      s603 <= s602;
      s604 <= s603;
      s605 <= s604;
      s606 <= s605;
      s607 <= s606;
      s608 <= s607;
      s609 <= s608;
      s610 <= s609;
      s611 <= s610;
      s612 <= s611;
      s613 <= s612;
      s614 <= s613;
      s615 <= s614;
      s616 <= s615;
      s617 <= s616;
      s618 <= s617;
      s619 <= s618;
      s620 <= s619;
      s621 <= s620;
      s622 <= s621;
      s623 <= s622;
      s624 <= s623;
      s625 <= s624;
      s626 <= s625;
      s627 <= s626;
      s628 <= s627;
      s629 <= s628;
      s630 <= s629;
      s631 <= s630;
      s632 <= s631;
      s633 <= s632;
      s634 <= s633;
      s635 <= s634;
      s636 <= s635;
      s637 <= s636;
      s638 <= s637;
      s639 <= s638;
      s640 <= s639;
      s641 <= s640;
      s642 <= s641;
      s643 <= s642;
      s644 <= s643;
      s645 <= s644;
      s646 <= s645;
      s647 <= s646;
      s648 <= s647;
      s649 <= s648;
      s650 <= s649;
      s651 <= s650;
      s652 <= s651;
      s653 <= s652;
      s654 <= s653;
      s655 <= s654;
      s656 <= s655;
      s657 <= s656;
      s658 <= s657;
      s659 <= s658;
      s660 <= s659;
      s661 <= s660;
      s662 <= s661;
      s663 <= s662;
      s664 <= s663;
      s665 <= s664;
      s666 <= s665;
      s667 <= s666;
      s668 <= s667;
      s669 <= s668;
      s670 <= s669;
      s671 <= s670;
      s672 <= s671;
      s673 <= s672;
      s674 <= s673;
      s675 <= s674;
      s676 <= s675;
      s677 <= s676;
      s678 <= s677;
      s679 <= s678;
      s680 <= s679;
      s681 <= s680;
      s682 <= s681;
      s683 <= s682;
      s684 <= s683;
      s685 <= s684;
      s686 <= s685;
      s687 <= s686;
      s688 <= s687;
      s689 <= s688;
      s690 <= s689;
      s691 <= s690;
      s692 <= s691;
      s693 <= s692;
      s694 <= s693;
      s695 <= s694;
      s696 <= s695;
      s697 <= s696;
      s698 <= s697;
      s699 <= s698;
      s700 <= s699;
      s701 <= s700;
      s702 <= s701;
      s703 <= s702;
      s704 <= s703;
      s705 <= s704;
      s706 <= s705;
      s707 <= s706;
      s708 <= s707;
      s709 <= s708;
      s710 <= s709;
      s711 <= s710;
      s712 <= s711;
      s713 <= s712;
      s714 <= s713;
      s715 <= s714;
      s716 <= s715;
      s717 <= s716;
      s718 <= s717;
      s719 <= s718;
      s720 <= s719;
      s721 <= s720;
      s722 <= s721;
      s723 <= s722;
      s724 <= s723;
      s725 <= s724;
      s726 <= s725;
      s727 <= s726;
      s728 <= s727;
      s729 <= s728;
      s730 <= s729;
      s731 <= s730;
      s732 <= s731;
      s733 <= s732;
      s734 <= s733;
      s735 <= s734;
      s736 <= s735;
      s737 <= s736;
      s738 <= s737;
      s739 <= s738;
      s740 <= s739;
      s741 <= s740;
      s742 <= s741;
      s743 <= s742;
      s744 <= s743;
      s745 <= s744;
      s746 <= s745;
      s747 <= s746;
      s748 <= s747;
      s749 <= s748;
      s750 <= s749;
      s751 <= s750;
      s752 <= s751;
      s753 <= s752;
      s754 <= s753;
      s755 <= s754;
      s756 <= s755;
      s757 <= s756;
      s758 <= s757;
      s759 <= s758;
      s760 <= s759;
      s761 <= s760;
      s762 <= s761;
      s763 <= s762;
      s764 <= s763;
      s765 <= s764;
      s766 <= s765;
      s767 <= s766;
      s768 <= s767;
      s769 <= s768;
      s770 <= s769;
      s771 <= s770;
      s772 <= s771;
      s773 <= s772;
      s774 <= s773;
      s775 <= s774;
      s776 <= s775;
      s777 <= s776;
      s778 <= s777;
      s779 <= s778;
      s780 <= s779;
      s781 <= s780;
      s782 <= s781;
      s783 <= s782;
      s784 <= s783;
      s785 <= s784;
      s786 <= s785;
      s787 <= s786;
      s788 <= s787;
      s789 <= s788;
      s790 <= s789;
      s791 <= s790;
      s792 <= s791;
      s793 <= s792;
      s794 <= s793;
      s795 <= s794;
      s796 <= s795;
      s797 <= s796;
      s798 <= s797;
      s799 <= s798;
      s800 <= s799;
      s801 <= s800;
      s802 <= s801;
      s803 <= s802;
      s804 <= s803;
      s805 <= s804;
      s806 <= s805;
      s807 <= s806;
      s808 <= s807;
      s809 <= s808;
      s810 <= s809;
      s811 <= s810;
      s812 <= s811;
      s813 <= s812;
      s814 <= s813;
      s815 <= s814;
      s816 <= s815;
      s817 <= s816;
      s818 <= s817;
      s819 <= s818;
      s820 <= s819;
      s821 <= s820;
      s822 <= s821;
      s823 <= s822;
      s824 <= s823;
      s825 <= s824;
      s826 <= s825;
      s827 <= s826;
      s828 <= s827;
      s829 <= s828;
      s830 <= s829;
      s831 <= s830;
      s832 <= s831;
      s833 <= s832;
      s834 <= s833;
      s835 <= s834;
      s836 <= s835;
      s837 <= s836;
      s838 <= s837;
      s839 <= s838;
      s840 <= s839;
      s841 <= s840;
      s842 <= s841;
      s843 <= s842;
      s844 <= s843;
      s845 <= s844;
      s846 <= s845;
      s847 <= s846;
      s848 <= s847;
      s849 <= s848;
      s850 <= s849;
      s851 <= s850;
      s852 <= s851;
      s853 <= s852;
      s854 <= s853;
      s855 <= s854;
      s856 <= s855;
      s857 <= s856;
      s858 <= s857;
      s859 <= s858;
      s860 <= s859;
      s861 <= s860;
      s862 <= s861;
      s863 <= s862;
      s864 <= s863;
      s865 <= s864;
      s866 <= s865;
      s867 <= s866;
      s868 <= s867;
      s869 <= s868;
      s870 <= s869;
      s871 <= s870;
      s872 <= s871;
      s873 <= s872;
      s874 <= s873;
      s875 <= s874;
      s876 <= s875;
      s877 <= s876;
      s878 <= s877;
      s879 <= s878;
      s880 <= s879;
      s881 <= s880;
      s882 <= s881;
      s883 <= s882;
      s884 <= s883;
      s885 <= s884;
      s886 <= s885;
      s887 <= s886;
      s888 <= s887;
      s889 <= s888;
      s890 <= s889;
      s891 <= s890;
      s892 <= s891;
      s893 <= s892;
      s894 <= s893;
      s895 <= s894;
      s896 <= s895;
      s897 <= s896;
      s898 <= s897;
      s899 <= s898;
      s900 <= s899;
      s901 <= s900;
      s902 <= s901;
      s903 <= s902;
      s904 <= s903;
      s905 <= s904;
      s906 <= s905;
      s907 <= s906;
      s908 <= s907;
      s909 <= s908;
      s910 <= s909;
      s911 <= s910;
      s912 <= s911;
      s913 <= s912;
      s914 <= s913;
      s915 <= s914;
      s916 <= s915;
      s917 <= s916;
      s918 <= s917;
      s919 <= s918;
      s920 <= s919;
      s921 <= s920;
      s922 <= s921;
      s923 <= s922;
      s924 <= s923;
      s925 <= s924;
      s926 <= s925;
      s927 <= s926;
      s928 <= s927;
      s929 <= s928;
      s930 <= s929;
      s931 <= s930;
      s932 <= s931;
      s933 <= s932;
      s934 <= s933;
      s935 <= s934;
      s936 <= s935;
      s937 <= s936;
      s938 <= s937;
      s939 <= s938;
      s940 <= s939;
      s941 <= s940;
      s942 <= s941;
      s943 <= s942;
      s944 <= s943;
      s945 <= s944;
      s946 <= s945;
      s947 <= s946;
      Y <= s947;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1016_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1016 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1016_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1016_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
signal s558 : std_logic_vector(33 downto 0) := (others => '0');
signal s559 : std_logic_vector(33 downto 0) := (others => '0');
signal s560 : std_logic_vector(33 downto 0) := (others => '0');
signal s561 : std_logic_vector(33 downto 0) := (others => '0');
signal s562 : std_logic_vector(33 downto 0) := (others => '0');
signal s563 : std_logic_vector(33 downto 0) := (others => '0');
signal s564 : std_logic_vector(33 downto 0) := (others => '0');
signal s565 : std_logic_vector(33 downto 0) := (others => '0');
signal s566 : std_logic_vector(33 downto 0) := (others => '0');
signal s567 : std_logic_vector(33 downto 0) := (others => '0');
signal s568 : std_logic_vector(33 downto 0) := (others => '0');
signal s569 : std_logic_vector(33 downto 0) := (others => '0');
signal s570 : std_logic_vector(33 downto 0) := (others => '0');
signal s571 : std_logic_vector(33 downto 0) := (others => '0');
signal s572 : std_logic_vector(33 downto 0) := (others => '0');
signal s573 : std_logic_vector(33 downto 0) := (others => '0');
signal s574 : std_logic_vector(33 downto 0) := (others => '0');
signal s575 : std_logic_vector(33 downto 0) := (others => '0');
signal s576 : std_logic_vector(33 downto 0) := (others => '0');
signal s577 : std_logic_vector(33 downto 0) := (others => '0');
signal s578 : std_logic_vector(33 downto 0) := (others => '0');
signal s579 : std_logic_vector(33 downto 0) := (others => '0');
signal s580 : std_logic_vector(33 downto 0) := (others => '0');
signal s581 : std_logic_vector(33 downto 0) := (others => '0');
signal s582 : std_logic_vector(33 downto 0) := (others => '0');
signal s583 : std_logic_vector(33 downto 0) := (others => '0');
signal s584 : std_logic_vector(33 downto 0) := (others => '0');
signal s585 : std_logic_vector(33 downto 0) := (others => '0');
signal s586 : std_logic_vector(33 downto 0) := (others => '0');
signal s587 : std_logic_vector(33 downto 0) := (others => '0');
signal s588 : std_logic_vector(33 downto 0) := (others => '0');
signal s589 : std_logic_vector(33 downto 0) := (others => '0');
signal s590 : std_logic_vector(33 downto 0) := (others => '0');
signal s591 : std_logic_vector(33 downto 0) := (others => '0');
signal s592 : std_logic_vector(33 downto 0) := (others => '0');
signal s593 : std_logic_vector(33 downto 0) := (others => '0');
signal s594 : std_logic_vector(33 downto 0) := (others => '0');
signal s595 : std_logic_vector(33 downto 0) := (others => '0');
signal s596 : std_logic_vector(33 downto 0) := (others => '0');
signal s597 : std_logic_vector(33 downto 0) := (others => '0');
signal s598 : std_logic_vector(33 downto 0) := (others => '0');
signal s599 : std_logic_vector(33 downto 0) := (others => '0');
signal s600 : std_logic_vector(33 downto 0) := (others => '0');
signal s601 : std_logic_vector(33 downto 0) := (others => '0');
signal s602 : std_logic_vector(33 downto 0) := (others => '0');
signal s603 : std_logic_vector(33 downto 0) := (others => '0');
signal s604 : std_logic_vector(33 downto 0) := (others => '0');
signal s605 : std_logic_vector(33 downto 0) := (others => '0');
signal s606 : std_logic_vector(33 downto 0) := (others => '0');
signal s607 : std_logic_vector(33 downto 0) := (others => '0');
signal s608 : std_logic_vector(33 downto 0) := (others => '0');
signal s609 : std_logic_vector(33 downto 0) := (others => '0');
signal s610 : std_logic_vector(33 downto 0) := (others => '0');
signal s611 : std_logic_vector(33 downto 0) := (others => '0');
signal s612 : std_logic_vector(33 downto 0) := (others => '0');
signal s613 : std_logic_vector(33 downto 0) := (others => '0');
signal s614 : std_logic_vector(33 downto 0) := (others => '0');
signal s615 : std_logic_vector(33 downto 0) := (others => '0');
signal s616 : std_logic_vector(33 downto 0) := (others => '0');
signal s617 : std_logic_vector(33 downto 0) := (others => '0');
signal s618 : std_logic_vector(33 downto 0) := (others => '0');
signal s619 : std_logic_vector(33 downto 0) := (others => '0');
signal s620 : std_logic_vector(33 downto 0) := (others => '0');
signal s621 : std_logic_vector(33 downto 0) := (others => '0');
signal s622 : std_logic_vector(33 downto 0) := (others => '0');
signal s623 : std_logic_vector(33 downto 0) := (others => '0');
signal s624 : std_logic_vector(33 downto 0) := (others => '0');
signal s625 : std_logic_vector(33 downto 0) := (others => '0');
signal s626 : std_logic_vector(33 downto 0) := (others => '0');
signal s627 : std_logic_vector(33 downto 0) := (others => '0');
signal s628 : std_logic_vector(33 downto 0) := (others => '0');
signal s629 : std_logic_vector(33 downto 0) := (others => '0');
signal s630 : std_logic_vector(33 downto 0) := (others => '0');
signal s631 : std_logic_vector(33 downto 0) := (others => '0');
signal s632 : std_logic_vector(33 downto 0) := (others => '0');
signal s633 : std_logic_vector(33 downto 0) := (others => '0');
signal s634 : std_logic_vector(33 downto 0) := (others => '0');
signal s635 : std_logic_vector(33 downto 0) := (others => '0');
signal s636 : std_logic_vector(33 downto 0) := (others => '0');
signal s637 : std_logic_vector(33 downto 0) := (others => '0');
signal s638 : std_logic_vector(33 downto 0) := (others => '0');
signal s639 : std_logic_vector(33 downto 0) := (others => '0');
signal s640 : std_logic_vector(33 downto 0) := (others => '0');
signal s641 : std_logic_vector(33 downto 0) := (others => '0');
signal s642 : std_logic_vector(33 downto 0) := (others => '0');
signal s643 : std_logic_vector(33 downto 0) := (others => '0');
signal s644 : std_logic_vector(33 downto 0) := (others => '0');
signal s645 : std_logic_vector(33 downto 0) := (others => '0');
signal s646 : std_logic_vector(33 downto 0) := (others => '0');
signal s647 : std_logic_vector(33 downto 0) := (others => '0');
signal s648 : std_logic_vector(33 downto 0) := (others => '0');
signal s649 : std_logic_vector(33 downto 0) := (others => '0');
signal s650 : std_logic_vector(33 downto 0) := (others => '0');
signal s651 : std_logic_vector(33 downto 0) := (others => '0');
signal s652 : std_logic_vector(33 downto 0) := (others => '0');
signal s653 : std_logic_vector(33 downto 0) := (others => '0');
signal s654 : std_logic_vector(33 downto 0) := (others => '0');
signal s655 : std_logic_vector(33 downto 0) := (others => '0');
signal s656 : std_logic_vector(33 downto 0) := (others => '0');
signal s657 : std_logic_vector(33 downto 0) := (others => '0');
signal s658 : std_logic_vector(33 downto 0) := (others => '0');
signal s659 : std_logic_vector(33 downto 0) := (others => '0');
signal s660 : std_logic_vector(33 downto 0) := (others => '0');
signal s661 : std_logic_vector(33 downto 0) := (others => '0');
signal s662 : std_logic_vector(33 downto 0) := (others => '0');
signal s663 : std_logic_vector(33 downto 0) := (others => '0');
signal s664 : std_logic_vector(33 downto 0) := (others => '0');
signal s665 : std_logic_vector(33 downto 0) := (others => '0');
signal s666 : std_logic_vector(33 downto 0) := (others => '0');
signal s667 : std_logic_vector(33 downto 0) := (others => '0');
signal s668 : std_logic_vector(33 downto 0) := (others => '0');
signal s669 : std_logic_vector(33 downto 0) := (others => '0');
signal s670 : std_logic_vector(33 downto 0) := (others => '0');
signal s671 : std_logic_vector(33 downto 0) := (others => '0');
signal s672 : std_logic_vector(33 downto 0) := (others => '0');
signal s673 : std_logic_vector(33 downto 0) := (others => '0');
signal s674 : std_logic_vector(33 downto 0) := (others => '0');
signal s675 : std_logic_vector(33 downto 0) := (others => '0');
signal s676 : std_logic_vector(33 downto 0) := (others => '0');
signal s677 : std_logic_vector(33 downto 0) := (others => '0');
signal s678 : std_logic_vector(33 downto 0) := (others => '0');
signal s679 : std_logic_vector(33 downto 0) := (others => '0');
signal s680 : std_logic_vector(33 downto 0) := (others => '0');
signal s681 : std_logic_vector(33 downto 0) := (others => '0');
signal s682 : std_logic_vector(33 downto 0) := (others => '0');
signal s683 : std_logic_vector(33 downto 0) := (others => '0');
signal s684 : std_logic_vector(33 downto 0) := (others => '0');
signal s685 : std_logic_vector(33 downto 0) := (others => '0');
signal s686 : std_logic_vector(33 downto 0) := (others => '0');
signal s687 : std_logic_vector(33 downto 0) := (others => '0');
signal s688 : std_logic_vector(33 downto 0) := (others => '0');
signal s689 : std_logic_vector(33 downto 0) := (others => '0');
signal s690 : std_logic_vector(33 downto 0) := (others => '0');
signal s691 : std_logic_vector(33 downto 0) := (others => '0');
signal s692 : std_logic_vector(33 downto 0) := (others => '0');
signal s693 : std_logic_vector(33 downto 0) := (others => '0');
signal s694 : std_logic_vector(33 downto 0) := (others => '0');
signal s695 : std_logic_vector(33 downto 0) := (others => '0');
signal s696 : std_logic_vector(33 downto 0) := (others => '0');
signal s697 : std_logic_vector(33 downto 0) := (others => '0');
signal s698 : std_logic_vector(33 downto 0) := (others => '0');
signal s699 : std_logic_vector(33 downto 0) := (others => '0');
signal s700 : std_logic_vector(33 downto 0) := (others => '0');
signal s701 : std_logic_vector(33 downto 0) := (others => '0');
signal s702 : std_logic_vector(33 downto 0) := (others => '0');
signal s703 : std_logic_vector(33 downto 0) := (others => '0');
signal s704 : std_logic_vector(33 downto 0) := (others => '0');
signal s705 : std_logic_vector(33 downto 0) := (others => '0');
signal s706 : std_logic_vector(33 downto 0) := (others => '0');
signal s707 : std_logic_vector(33 downto 0) := (others => '0');
signal s708 : std_logic_vector(33 downto 0) := (others => '0');
signal s709 : std_logic_vector(33 downto 0) := (others => '0');
signal s710 : std_logic_vector(33 downto 0) := (others => '0');
signal s711 : std_logic_vector(33 downto 0) := (others => '0');
signal s712 : std_logic_vector(33 downto 0) := (others => '0');
signal s713 : std_logic_vector(33 downto 0) := (others => '0');
signal s714 : std_logic_vector(33 downto 0) := (others => '0');
signal s715 : std_logic_vector(33 downto 0) := (others => '0');
signal s716 : std_logic_vector(33 downto 0) := (others => '0');
signal s717 : std_logic_vector(33 downto 0) := (others => '0');
signal s718 : std_logic_vector(33 downto 0) := (others => '0');
signal s719 : std_logic_vector(33 downto 0) := (others => '0');
signal s720 : std_logic_vector(33 downto 0) := (others => '0');
signal s721 : std_logic_vector(33 downto 0) := (others => '0');
signal s722 : std_logic_vector(33 downto 0) := (others => '0');
signal s723 : std_logic_vector(33 downto 0) := (others => '0');
signal s724 : std_logic_vector(33 downto 0) := (others => '0');
signal s725 : std_logic_vector(33 downto 0) := (others => '0');
signal s726 : std_logic_vector(33 downto 0) := (others => '0');
signal s727 : std_logic_vector(33 downto 0) := (others => '0');
signal s728 : std_logic_vector(33 downto 0) := (others => '0');
signal s729 : std_logic_vector(33 downto 0) := (others => '0');
signal s730 : std_logic_vector(33 downto 0) := (others => '0');
signal s731 : std_logic_vector(33 downto 0) := (others => '0');
signal s732 : std_logic_vector(33 downto 0) := (others => '0');
signal s733 : std_logic_vector(33 downto 0) := (others => '0');
signal s734 : std_logic_vector(33 downto 0) := (others => '0');
signal s735 : std_logic_vector(33 downto 0) := (others => '0');
signal s736 : std_logic_vector(33 downto 0) := (others => '0');
signal s737 : std_logic_vector(33 downto 0) := (others => '0');
signal s738 : std_logic_vector(33 downto 0) := (others => '0');
signal s739 : std_logic_vector(33 downto 0) := (others => '0');
signal s740 : std_logic_vector(33 downto 0) := (others => '0');
signal s741 : std_logic_vector(33 downto 0) := (others => '0');
signal s742 : std_logic_vector(33 downto 0) := (others => '0');
signal s743 : std_logic_vector(33 downto 0) := (others => '0');
signal s744 : std_logic_vector(33 downto 0) := (others => '0');
signal s745 : std_logic_vector(33 downto 0) := (others => '0');
signal s746 : std_logic_vector(33 downto 0) := (others => '0');
signal s747 : std_logic_vector(33 downto 0) := (others => '0');
signal s748 : std_logic_vector(33 downto 0) := (others => '0');
signal s749 : std_logic_vector(33 downto 0) := (others => '0');
signal s750 : std_logic_vector(33 downto 0) := (others => '0');
signal s751 : std_logic_vector(33 downto 0) := (others => '0');
signal s752 : std_logic_vector(33 downto 0) := (others => '0');
signal s753 : std_logic_vector(33 downto 0) := (others => '0');
signal s754 : std_logic_vector(33 downto 0) := (others => '0');
signal s755 : std_logic_vector(33 downto 0) := (others => '0');
signal s756 : std_logic_vector(33 downto 0) := (others => '0');
signal s757 : std_logic_vector(33 downto 0) := (others => '0');
signal s758 : std_logic_vector(33 downto 0) := (others => '0');
signal s759 : std_logic_vector(33 downto 0) := (others => '0');
signal s760 : std_logic_vector(33 downto 0) := (others => '0');
signal s761 : std_logic_vector(33 downto 0) := (others => '0');
signal s762 : std_logic_vector(33 downto 0) := (others => '0');
signal s763 : std_logic_vector(33 downto 0) := (others => '0');
signal s764 : std_logic_vector(33 downto 0) := (others => '0');
signal s765 : std_logic_vector(33 downto 0) := (others => '0');
signal s766 : std_logic_vector(33 downto 0) := (others => '0');
signal s767 : std_logic_vector(33 downto 0) := (others => '0');
signal s768 : std_logic_vector(33 downto 0) := (others => '0');
signal s769 : std_logic_vector(33 downto 0) := (others => '0');
signal s770 : std_logic_vector(33 downto 0) := (others => '0');
signal s771 : std_logic_vector(33 downto 0) := (others => '0');
signal s772 : std_logic_vector(33 downto 0) := (others => '0');
signal s773 : std_logic_vector(33 downto 0) := (others => '0');
signal s774 : std_logic_vector(33 downto 0) := (others => '0');
signal s775 : std_logic_vector(33 downto 0) := (others => '0');
signal s776 : std_logic_vector(33 downto 0) := (others => '0');
signal s777 : std_logic_vector(33 downto 0) := (others => '0');
signal s778 : std_logic_vector(33 downto 0) := (others => '0');
signal s779 : std_logic_vector(33 downto 0) := (others => '0');
signal s780 : std_logic_vector(33 downto 0) := (others => '0');
signal s781 : std_logic_vector(33 downto 0) := (others => '0');
signal s782 : std_logic_vector(33 downto 0) := (others => '0');
signal s783 : std_logic_vector(33 downto 0) := (others => '0');
signal s784 : std_logic_vector(33 downto 0) := (others => '0');
signal s785 : std_logic_vector(33 downto 0) := (others => '0');
signal s786 : std_logic_vector(33 downto 0) := (others => '0');
signal s787 : std_logic_vector(33 downto 0) := (others => '0');
signal s788 : std_logic_vector(33 downto 0) := (others => '0');
signal s789 : std_logic_vector(33 downto 0) := (others => '0');
signal s790 : std_logic_vector(33 downto 0) := (others => '0');
signal s791 : std_logic_vector(33 downto 0) := (others => '0');
signal s792 : std_logic_vector(33 downto 0) := (others => '0');
signal s793 : std_logic_vector(33 downto 0) := (others => '0');
signal s794 : std_logic_vector(33 downto 0) := (others => '0');
signal s795 : std_logic_vector(33 downto 0) := (others => '0');
signal s796 : std_logic_vector(33 downto 0) := (others => '0');
signal s797 : std_logic_vector(33 downto 0) := (others => '0');
signal s798 : std_logic_vector(33 downto 0) := (others => '0');
signal s799 : std_logic_vector(33 downto 0) := (others => '0');
signal s800 : std_logic_vector(33 downto 0) := (others => '0');
signal s801 : std_logic_vector(33 downto 0) := (others => '0');
signal s802 : std_logic_vector(33 downto 0) := (others => '0');
signal s803 : std_logic_vector(33 downto 0) := (others => '0');
signal s804 : std_logic_vector(33 downto 0) := (others => '0');
signal s805 : std_logic_vector(33 downto 0) := (others => '0');
signal s806 : std_logic_vector(33 downto 0) := (others => '0');
signal s807 : std_logic_vector(33 downto 0) := (others => '0');
signal s808 : std_logic_vector(33 downto 0) := (others => '0');
signal s809 : std_logic_vector(33 downto 0) := (others => '0');
signal s810 : std_logic_vector(33 downto 0) := (others => '0');
signal s811 : std_logic_vector(33 downto 0) := (others => '0');
signal s812 : std_logic_vector(33 downto 0) := (others => '0');
signal s813 : std_logic_vector(33 downto 0) := (others => '0');
signal s814 : std_logic_vector(33 downto 0) := (others => '0');
signal s815 : std_logic_vector(33 downto 0) := (others => '0');
signal s816 : std_logic_vector(33 downto 0) := (others => '0');
signal s817 : std_logic_vector(33 downto 0) := (others => '0');
signal s818 : std_logic_vector(33 downto 0) := (others => '0');
signal s819 : std_logic_vector(33 downto 0) := (others => '0');
signal s820 : std_logic_vector(33 downto 0) := (others => '0');
signal s821 : std_logic_vector(33 downto 0) := (others => '0');
signal s822 : std_logic_vector(33 downto 0) := (others => '0');
signal s823 : std_logic_vector(33 downto 0) := (others => '0');
signal s824 : std_logic_vector(33 downto 0) := (others => '0');
signal s825 : std_logic_vector(33 downto 0) := (others => '0');
signal s826 : std_logic_vector(33 downto 0) := (others => '0');
signal s827 : std_logic_vector(33 downto 0) := (others => '0');
signal s828 : std_logic_vector(33 downto 0) := (others => '0');
signal s829 : std_logic_vector(33 downto 0) := (others => '0');
signal s830 : std_logic_vector(33 downto 0) := (others => '0');
signal s831 : std_logic_vector(33 downto 0) := (others => '0');
signal s832 : std_logic_vector(33 downto 0) := (others => '0');
signal s833 : std_logic_vector(33 downto 0) := (others => '0');
signal s834 : std_logic_vector(33 downto 0) := (others => '0');
signal s835 : std_logic_vector(33 downto 0) := (others => '0');
signal s836 : std_logic_vector(33 downto 0) := (others => '0');
signal s837 : std_logic_vector(33 downto 0) := (others => '0');
signal s838 : std_logic_vector(33 downto 0) := (others => '0');
signal s839 : std_logic_vector(33 downto 0) := (others => '0');
signal s840 : std_logic_vector(33 downto 0) := (others => '0');
signal s841 : std_logic_vector(33 downto 0) := (others => '0');
signal s842 : std_logic_vector(33 downto 0) := (others => '0');
signal s843 : std_logic_vector(33 downto 0) := (others => '0');
signal s844 : std_logic_vector(33 downto 0) := (others => '0');
signal s845 : std_logic_vector(33 downto 0) := (others => '0');
signal s846 : std_logic_vector(33 downto 0) := (others => '0');
signal s847 : std_logic_vector(33 downto 0) := (others => '0');
signal s848 : std_logic_vector(33 downto 0) := (others => '0');
signal s849 : std_logic_vector(33 downto 0) := (others => '0');
signal s850 : std_logic_vector(33 downto 0) := (others => '0');
signal s851 : std_logic_vector(33 downto 0) := (others => '0');
signal s852 : std_logic_vector(33 downto 0) := (others => '0');
signal s853 : std_logic_vector(33 downto 0) := (others => '0');
signal s854 : std_logic_vector(33 downto 0) := (others => '0');
signal s855 : std_logic_vector(33 downto 0) := (others => '0');
signal s856 : std_logic_vector(33 downto 0) := (others => '0');
signal s857 : std_logic_vector(33 downto 0) := (others => '0');
signal s858 : std_logic_vector(33 downto 0) := (others => '0');
signal s859 : std_logic_vector(33 downto 0) := (others => '0');
signal s860 : std_logic_vector(33 downto 0) := (others => '0');
signal s861 : std_logic_vector(33 downto 0) := (others => '0');
signal s862 : std_logic_vector(33 downto 0) := (others => '0');
signal s863 : std_logic_vector(33 downto 0) := (others => '0');
signal s864 : std_logic_vector(33 downto 0) := (others => '0');
signal s865 : std_logic_vector(33 downto 0) := (others => '0');
signal s866 : std_logic_vector(33 downto 0) := (others => '0');
signal s867 : std_logic_vector(33 downto 0) := (others => '0');
signal s868 : std_logic_vector(33 downto 0) := (others => '0');
signal s869 : std_logic_vector(33 downto 0) := (others => '0');
signal s870 : std_logic_vector(33 downto 0) := (others => '0');
signal s871 : std_logic_vector(33 downto 0) := (others => '0');
signal s872 : std_logic_vector(33 downto 0) := (others => '0');
signal s873 : std_logic_vector(33 downto 0) := (others => '0');
signal s874 : std_logic_vector(33 downto 0) := (others => '0');
signal s875 : std_logic_vector(33 downto 0) := (others => '0');
signal s876 : std_logic_vector(33 downto 0) := (others => '0');
signal s877 : std_logic_vector(33 downto 0) := (others => '0');
signal s878 : std_logic_vector(33 downto 0) := (others => '0');
signal s879 : std_logic_vector(33 downto 0) := (others => '0');
signal s880 : std_logic_vector(33 downto 0) := (others => '0');
signal s881 : std_logic_vector(33 downto 0) := (others => '0');
signal s882 : std_logic_vector(33 downto 0) := (others => '0');
signal s883 : std_logic_vector(33 downto 0) := (others => '0');
signal s884 : std_logic_vector(33 downto 0) := (others => '0');
signal s885 : std_logic_vector(33 downto 0) := (others => '0');
signal s886 : std_logic_vector(33 downto 0) := (others => '0');
signal s887 : std_logic_vector(33 downto 0) := (others => '0');
signal s888 : std_logic_vector(33 downto 0) := (others => '0');
signal s889 : std_logic_vector(33 downto 0) := (others => '0');
signal s890 : std_logic_vector(33 downto 0) := (others => '0');
signal s891 : std_logic_vector(33 downto 0) := (others => '0');
signal s892 : std_logic_vector(33 downto 0) := (others => '0');
signal s893 : std_logic_vector(33 downto 0) := (others => '0');
signal s894 : std_logic_vector(33 downto 0) := (others => '0');
signal s895 : std_logic_vector(33 downto 0) := (others => '0');
signal s896 : std_logic_vector(33 downto 0) := (others => '0');
signal s897 : std_logic_vector(33 downto 0) := (others => '0');
signal s898 : std_logic_vector(33 downto 0) := (others => '0');
signal s899 : std_logic_vector(33 downto 0) := (others => '0');
signal s900 : std_logic_vector(33 downto 0) := (others => '0');
signal s901 : std_logic_vector(33 downto 0) := (others => '0');
signal s902 : std_logic_vector(33 downto 0) := (others => '0');
signal s903 : std_logic_vector(33 downto 0) := (others => '0');
signal s904 : std_logic_vector(33 downto 0) := (others => '0');
signal s905 : std_logic_vector(33 downto 0) := (others => '0');
signal s906 : std_logic_vector(33 downto 0) := (others => '0');
signal s907 : std_logic_vector(33 downto 0) := (others => '0');
signal s908 : std_logic_vector(33 downto 0) := (others => '0');
signal s909 : std_logic_vector(33 downto 0) := (others => '0');
signal s910 : std_logic_vector(33 downto 0) := (others => '0');
signal s911 : std_logic_vector(33 downto 0) := (others => '0');
signal s912 : std_logic_vector(33 downto 0) := (others => '0');
signal s913 : std_logic_vector(33 downto 0) := (others => '0');
signal s914 : std_logic_vector(33 downto 0) := (others => '0');
signal s915 : std_logic_vector(33 downto 0) := (others => '0');
signal s916 : std_logic_vector(33 downto 0) := (others => '0');
signal s917 : std_logic_vector(33 downto 0) := (others => '0');
signal s918 : std_logic_vector(33 downto 0) := (others => '0');
signal s919 : std_logic_vector(33 downto 0) := (others => '0');
signal s920 : std_logic_vector(33 downto 0) := (others => '0');
signal s921 : std_logic_vector(33 downto 0) := (others => '0');
signal s922 : std_logic_vector(33 downto 0) := (others => '0');
signal s923 : std_logic_vector(33 downto 0) := (others => '0');
signal s924 : std_logic_vector(33 downto 0) := (others => '0');
signal s925 : std_logic_vector(33 downto 0) := (others => '0');
signal s926 : std_logic_vector(33 downto 0) := (others => '0');
signal s927 : std_logic_vector(33 downto 0) := (others => '0');
signal s928 : std_logic_vector(33 downto 0) := (others => '0');
signal s929 : std_logic_vector(33 downto 0) := (others => '0');
signal s930 : std_logic_vector(33 downto 0) := (others => '0');
signal s931 : std_logic_vector(33 downto 0) := (others => '0');
signal s932 : std_logic_vector(33 downto 0) := (others => '0');
signal s933 : std_logic_vector(33 downto 0) := (others => '0');
signal s934 : std_logic_vector(33 downto 0) := (others => '0');
signal s935 : std_logic_vector(33 downto 0) := (others => '0');
signal s936 : std_logic_vector(33 downto 0) := (others => '0');
signal s937 : std_logic_vector(33 downto 0) := (others => '0');
signal s938 : std_logic_vector(33 downto 0) := (others => '0');
signal s939 : std_logic_vector(33 downto 0) := (others => '0');
signal s940 : std_logic_vector(33 downto 0) := (others => '0');
signal s941 : std_logic_vector(33 downto 0) := (others => '0');
signal s942 : std_logic_vector(33 downto 0) := (others => '0');
signal s943 : std_logic_vector(33 downto 0) := (others => '0');
signal s944 : std_logic_vector(33 downto 0) := (others => '0');
signal s945 : std_logic_vector(33 downto 0) := (others => '0');
signal s946 : std_logic_vector(33 downto 0) := (others => '0');
signal s947 : std_logic_vector(33 downto 0) := (others => '0');
signal s948 : std_logic_vector(33 downto 0) := (others => '0');
signal s949 : std_logic_vector(33 downto 0) := (others => '0');
signal s950 : std_logic_vector(33 downto 0) := (others => '0');
signal s951 : std_logic_vector(33 downto 0) := (others => '0');
signal s952 : std_logic_vector(33 downto 0) := (others => '0');
signal s953 : std_logic_vector(33 downto 0) := (others => '0');
signal s954 : std_logic_vector(33 downto 0) := (others => '0');
signal s955 : std_logic_vector(33 downto 0) := (others => '0');
signal s956 : std_logic_vector(33 downto 0) := (others => '0');
signal s957 : std_logic_vector(33 downto 0) := (others => '0');
signal s958 : std_logic_vector(33 downto 0) := (others => '0');
signal s959 : std_logic_vector(33 downto 0) := (others => '0');
signal s960 : std_logic_vector(33 downto 0) := (others => '0');
signal s961 : std_logic_vector(33 downto 0) := (others => '0');
signal s962 : std_logic_vector(33 downto 0) := (others => '0');
signal s963 : std_logic_vector(33 downto 0) := (others => '0');
signal s964 : std_logic_vector(33 downto 0) := (others => '0');
signal s965 : std_logic_vector(33 downto 0) := (others => '0');
signal s966 : std_logic_vector(33 downto 0) := (others => '0');
signal s967 : std_logic_vector(33 downto 0) := (others => '0');
signal s968 : std_logic_vector(33 downto 0) := (others => '0');
signal s969 : std_logic_vector(33 downto 0) := (others => '0');
signal s970 : std_logic_vector(33 downto 0) := (others => '0');
signal s971 : std_logic_vector(33 downto 0) := (others => '0');
signal s972 : std_logic_vector(33 downto 0) := (others => '0');
signal s973 : std_logic_vector(33 downto 0) := (others => '0');
signal s974 : std_logic_vector(33 downto 0) := (others => '0');
signal s975 : std_logic_vector(33 downto 0) := (others => '0');
signal s976 : std_logic_vector(33 downto 0) := (others => '0');
signal s977 : std_logic_vector(33 downto 0) := (others => '0');
signal s978 : std_logic_vector(33 downto 0) := (others => '0');
signal s979 : std_logic_vector(33 downto 0) := (others => '0');
signal s980 : std_logic_vector(33 downto 0) := (others => '0');
signal s981 : std_logic_vector(33 downto 0) := (others => '0');
signal s982 : std_logic_vector(33 downto 0) := (others => '0');
signal s983 : std_logic_vector(33 downto 0) := (others => '0');
signal s984 : std_logic_vector(33 downto 0) := (others => '0');
signal s985 : std_logic_vector(33 downto 0) := (others => '0');
signal s986 : std_logic_vector(33 downto 0) := (others => '0');
signal s987 : std_logic_vector(33 downto 0) := (others => '0');
signal s988 : std_logic_vector(33 downto 0) := (others => '0');
signal s989 : std_logic_vector(33 downto 0) := (others => '0');
signal s990 : std_logic_vector(33 downto 0) := (others => '0');
signal s991 : std_logic_vector(33 downto 0) := (others => '0');
signal s992 : std_logic_vector(33 downto 0) := (others => '0');
signal s993 : std_logic_vector(33 downto 0) := (others => '0');
signal s994 : std_logic_vector(33 downto 0) := (others => '0');
signal s995 : std_logic_vector(33 downto 0) := (others => '0');
signal s996 : std_logic_vector(33 downto 0) := (others => '0');
signal s997 : std_logic_vector(33 downto 0) := (others => '0');
signal s998 : std_logic_vector(33 downto 0) := (others => '0');
signal s999 : std_logic_vector(33 downto 0) := (others => '0');
signal s1000 : std_logic_vector(33 downto 0) := (others => '0');
signal s1001 : std_logic_vector(33 downto 0) := (others => '0');
signal s1002 : std_logic_vector(33 downto 0) := (others => '0');
signal s1003 : std_logic_vector(33 downto 0) := (others => '0');
signal s1004 : std_logic_vector(33 downto 0) := (others => '0');
signal s1005 : std_logic_vector(33 downto 0) := (others => '0');
signal s1006 : std_logic_vector(33 downto 0) := (others => '0');
signal s1007 : std_logic_vector(33 downto 0) := (others => '0');
signal s1008 : std_logic_vector(33 downto 0) := (others => '0');
signal s1009 : std_logic_vector(33 downto 0) := (others => '0');
signal s1010 : std_logic_vector(33 downto 0) := (others => '0');
signal s1011 : std_logic_vector(33 downto 0) := (others => '0');
signal s1012 : std_logic_vector(33 downto 0) := (others => '0');
signal s1013 : std_logic_vector(33 downto 0) := (others => '0');
signal s1014 : std_logic_vector(33 downto 0) := (others => '0');
signal s1015 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
      s558 <= "0000000000000000000000000000000000";
      s559 <= "0000000000000000000000000000000000";
      s560 <= "0000000000000000000000000000000000";
      s561 <= "0000000000000000000000000000000000";
      s562 <= "0000000000000000000000000000000000";
      s563 <= "0000000000000000000000000000000000";
      s564 <= "0000000000000000000000000000000000";
      s565 <= "0000000000000000000000000000000000";
      s566 <= "0000000000000000000000000000000000";
      s567 <= "0000000000000000000000000000000000";
      s568 <= "0000000000000000000000000000000000";
      s569 <= "0000000000000000000000000000000000";
      s570 <= "0000000000000000000000000000000000";
      s571 <= "0000000000000000000000000000000000";
      s572 <= "0000000000000000000000000000000000";
      s573 <= "0000000000000000000000000000000000";
      s574 <= "0000000000000000000000000000000000";
      s575 <= "0000000000000000000000000000000000";
      s576 <= "0000000000000000000000000000000000";
      s577 <= "0000000000000000000000000000000000";
      s578 <= "0000000000000000000000000000000000";
      s579 <= "0000000000000000000000000000000000";
      s580 <= "0000000000000000000000000000000000";
      s581 <= "0000000000000000000000000000000000";
      s582 <= "0000000000000000000000000000000000";
      s583 <= "0000000000000000000000000000000000";
      s584 <= "0000000000000000000000000000000000";
      s585 <= "0000000000000000000000000000000000";
      s586 <= "0000000000000000000000000000000000";
      s587 <= "0000000000000000000000000000000000";
      s588 <= "0000000000000000000000000000000000";
      s589 <= "0000000000000000000000000000000000";
      s590 <= "0000000000000000000000000000000000";
      s591 <= "0000000000000000000000000000000000";
      s592 <= "0000000000000000000000000000000000";
      s593 <= "0000000000000000000000000000000000";
      s594 <= "0000000000000000000000000000000000";
      s595 <= "0000000000000000000000000000000000";
      s596 <= "0000000000000000000000000000000000";
      s597 <= "0000000000000000000000000000000000";
      s598 <= "0000000000000000000000000000000000";
      s599 <= "0000000000000000000000000000000000";
      s600 <= "0000000000000000000000000000000000";
      s601 <= "0000000000000000000000000000000000";
      s602 <= "0000000000000000000000000000000000";
      s603 <= "0000000000000000000000000000000000";
      s604 <= "0000000000000000000000000000000000";
      s605 <= "0000000000000000000000000000000000";
      s606 <= "0000000000000000000000000000000000";
      s607 <= "0000000000000000000000000000000000";
      s608 <= "0000000000000000000000000000000000";
      s609 <= "0000000000000000000000000000000000";
      s610 <= "0000000000000000000000000000000000";
      s611 <= "0000000000000000000000000000000000";
      s612 <= "0000000000000000000000000000000000";
      s613 <= "0000000000000000000000000000000000";
      s614 <= "0000000000000000000000000000000000";
      s615 <= "0000000000000000000000000000000000";
      s616 <= "0000000000000000000000000000000000";
      s617 <= "0000000000000000000000000000000000";
      s618 <= "0000000000000000000000000000000000";
      s619 <= "0000000000000000000000000000000000";
      s620 <= "0000000000000000000000000000000000";
      s621 <= "0000000000000000000000000000000000";
      s622 <= "0000000000000000000000000000000000";
      s623 <= "0000000000000000000000000000000000";
      s624 <= "0000000000000000000000000000000000";
      s625 <= "0000000000000000000000000000000000";
      s626 <= "0000000000000000000000000000000000";
      s627 <= "0000000000000000000000000000000000";
      s628 <= "0000000000000000000000000000000000";
      s629 <= "0000000000000000000000000000000000";
      s630 <= "0000000000000000000000000000000000";
      s631 <= "0000000000000000000000000000000000";
      s632 <= "0000000000000000000000000000000000";
      s633 <= "0000000000000000000000000000000000";
      s634 <= "0000000000000000000000000000000000";
      s635 <= "0000000000000000000000000000000000";
      s636 <= "0000000000000000000000000000000000";
      s637 <= "0000000000000000000000000000000000";
      s638 <= "0000000000000000000000000000000000";
      s639 <= "0000000000000000000000000000000000";
      s640 <= "0000000000000000000000000000000000";
      s641 <= "0000000000000000000000000000000000";
      s642 <= "0000000000000000000000000000000000";
      s643 <= "0000000000000000000000000000000000";
      s644 <= "0000000000000000000000000000000000";
      s645 <= "0000000000000000000000000000000000";
      s646 <= "0000000000000000000000000000000000";
      s647 <= "0000000000000000000000000000000000";
      s648 <= "0000000000000000000000000000000000";
      s649 <= "0000000000000000000000000000000000";
      s650 <= "0000000000000000000000000000000000";
      s651 <= "0000000000000000000000000000000000";
      s652 <= "0000000000000000000000000000000000";
      s653 <= "0000000000000000000000000000000000";
      s654 <= "0000000000000000000000000000000000";
      s655 <= "0000000000000000000000000000000000";
      s656 <= "0000000000000000000000000000000000";
      s657 <= "0000000000000000000000000000000000";
      s658 <= "0000000000000000000000000000000000";
      s659 <= "0000000000000000000000000000000000";
      s660 <= "0000000000000000000000000000000000";
      s661 <= "0000000000000000000000000000000000";
      s662 <= "0000000000000000000000000000000000";
      s663 <= "0000000000000000000000000000000000";
      s664 <= "0000000000000000000000000000000000";
      s665 <= "0000000000000000000000000000000000";
      s666 <= "0000000000000000000000000000000000";
      s667 <= "0000000000000000000000000000000000";
      s668 <= "0000000000000000000000000000000000";
      s669 <= "0000000000000000000000000000000000";
      s670 <= "0000000000000000000000000000000000";
      s671 <= "0000000000000000000000000000000000";
      s672 <= "0000000000000000000000000000000000";
      s673 <= "0000000000000000000000000000000000";
      s674 <= "0000000000000000000000000000000000";
      s675 <= "0000000000000000000000000000000000";
      s676 <= "0000000000000000000000000000000000";
      s677 <= "0000000000000000000000000000000000";
      s678 <= "0000000000000000000000000000000000";
      s679 <= "0000000000000000000000000000000000";
      s680 <= "0000000000000000000000000000000000";
      s681 <= "0000000000000000000000000000000000";
      s682 <= "0000000000000000000000000000000000";
      s683 <= "0000000000000000000000000000000000";
      s684 <= "0000000000000000000000000000000000";
      s685 <= "0000000000000000000000000000000000";
      s686 <= "0000000000000000000000000000000000";
      s687 <= "0000000000000000000000000000000000";
      s688 <= "0000000000000000000000000000000000";
      s689 <= "0000000000000000000000000000000000";
      s690 <= "0000000000000000000000000000000000";
      s691 <= "0000000000000000000000000000000000";
      s692 <= "0000000000000000000000000000000000";
      s693 <= "0000000000000000000000000000000000";
      s694 <= "0000000000000000000000000000000000";
      s695 <= "0000000000000000000000000000000000";
      s696 <= "0000000000000000000000000000000000";
      s697 <= "0000000000000000000000000000000000";
      s698 <= "0000000000000000000000000000000000";
      s699 <= "0000000000000000000000000000000000";
      s700 <= "0000000000000000000000000000000000";
      s701 <= "0000000000000000000000000000000000";
      s702 <= "0000000000000000000000000000000000";
      s703 <= "0000000000000000000000000000000000";
      s704 <= "0000000000000000000000000000000000";
      s705 <= "0000000000000000000000000000000000";
      s706 <= "0000000000000000000000000000000000";
      s707 <= "0000000000000000000000000000000000";
      s708 <= "0000000000000000000000000000000000";
      s709 <= "0000000000000000000000000000000000";
      s710 <= "0000000000000000000000000000000000";
      s711 <= "0000000000000000000000000000000000";
      s712 <= "0000000000000000000000000000000000";
      s713 <= "0000000000000000000000000000000000";
      s714 <= "0000000000000000000000000000000000";
      s715 <= "0000000000000000000000000000000000";
      s716 <= "0000000000000000000000000000000000";
      s717 <= "0000000000000000000000000000000000";
      s718 <= "0000000000000000000000000000000000";
      s719 <= "0000000000000000000000000000000000";
      s720 <= "0000000000000000000000000000000000";
      s721 <= "0000000000000000000000000000000000";
      s722 <= "0000000000000000000000000000000000";
      s723 <= "0000000000000000000000000000000000";
      s724 <= "0000000000000000000000000000000000";
      s725 <= "0000000000000000000000000000000000";
      s726 <= "0000000000000000000000000000000000";
      s727 <= "0000000000000000000000000000000000";
      s728 <= "0000000000000000000000000000000000";
      s729 <= "0000000000000000000000000000000000";
      s730 <= "0000000000000000000000000000000000";
      s731 <= "0000000000000000000000000000000000";
      s732 <= "0000000000000000000000000000000000";
      s733 <= "0000000000000000000000000000000000";
      s734 <= "0000000000000000000000000000000000";
      s735 <= "0000000000000000000000000000000000";
      s736 <= "0000000000000000000000000000000000";
      s737 <= "0000000000000000000000000000000000";
      s738 <= "0000000000000000000000000000000000";
      s739 <= "0000000000000000000000000000000000";
      s740 <= "0000000000000000000000000000000000";
      s741 <= "0000000000000000000000000000000000";
      s742 <= "0000000000000000000000000000000000";
      s743 <= "0000000000000000000000000000000000";
      s744 <= "0000000000000000000000000000000000";
      s745 <= "0000000000000000000000000000000000";
      s746 <= "0000000000000000000000000000000000";
      s747 <= "0000000000000000000000000000000000";
      s748 <= "0000000000000000000000000000000000";
      s749 <= "0000000000000000000000000000000000";
      s750 <= "0000000000000000000000000000000000";
      s751 <= "0000000000000000000000000000000000";
      s752 <= "0000000000000000000000000000000000";
      s753 <= "0000000000000000000000000000000000";
      s754 <= "0000000000000000000000000000000000";
      s755 <= "0000000000000000000000000000000000";
      s756 <= "0000000000000000000000000000000000";
      s757 <= "0000000000000000000000000000000000";
      s758 <= "0000000000000000000000000000000000";
      s759 <= "0000000000000000000000000000000000";
      s760 <= "0000000000000000000000000000000000";
      s761 <= "0000000000000000000000000000000000";
      s762 <= "0000000000000000000000000000000000";
      s763 <= "0000000000000000000000000000000000";
      s764 <= "0000000000000000000000000000000000";
      s765 <= "0000000000000000000000000000000000";
      s766 <= "0000000000000000000000000000000000";
      s767 <= "0000000000000000000000000000000000";
      s768 <= "0000000000000000000000000000000000";
      s769 <= "0000000000000000000000000000000000";
      s770 <= "0000000000000000000000000000000000";
      s771 <= "0000000000000000000000000000000000";
      s772 <= "0000000000000000000000000000000000";
      s773 <= "0000000000000000000000000000000000";
      s774 <= "0000000000000000000000000000000000";
      s775 <= "0000000000000000000000000000000000";
      s776 <= "0000000000000000000000000000000000";
      s777 <= "0000000000000000000000000000000000";
      s778 <= "0000000000000000000000000000000000";
      s779 <= "0000000000000000000000000000000000";
      s780 <= "0000000000000000000000000000000000";
      s781 <= "0000000000000000000000000000000000";
      s782 <= "0000000000000000000000000000000000";
      s783 <= "0000000000000000000000000000000000";
      s784 <= "0000000000000000000000000000000000";
      s785 <= "0000000000000000000000000000000000";
      s786 <= "0000000000000000000000000000000000";
      s787 <= "0000000000000000000000000000000000";
      s788 <= "0000000000000000000000000000000000";
      s789 <= "0000000000000000000000000000000000";
      s790 <= "0000000000000000000000000000000000";
      s791 <= "0000000000000000000000000000000000";
      s792 <= "0000000000000000000000000000000000";
      s793 <= "0000000000000000000000000000000000";
      s794 <= "0000000000000000000000000000000000";
      s795 <= "0000000000000000000000000000000000";
      s796 <= "0000000000000000000000000000000000";
      s797 <= "0000000000000000000000000000000000";
      s798 <= "0000000000000000000000000000000000";
      s799 <= "0000000000000000000000000000000000";
      s800 <= "0000000000000000000000000000000000";
      s801 <= "0000000000000000000000000000000000";
      s802 <= "0000000000000000000000000000000000";
      s803 <= "0000000000000000000000000000000000";
      s804 <= "0000000000000000000000000000000000";
      s805 <= "0000000000000000000000000000000000";
      s806 <= "0000000000000000000000000000000000";
      s807 <= "0000000000000000000000000000000000";
      s808 <= "0000000000000000000000000000000000";
      s809 <= "0000000000000000000000000000000000";
      s810 <= "0000000000000000000000000000000000";
      s811 <= "0000000000000000000000000000000000";
      s812 <= "0000000000000000000000000000000000";
      s813 <= "0000000000000000000000000000000000";
      s814 <= "0000000000000000000000000000000000";
      s815 <= "0000000000000000000000000000000000";
      s816 <= "0000000000000000000000000000000000";
      s817 <= "0000000000000000000000000000000000";
      s818 <= "0000000000000000000000000000000000";
      s819 <= "0000000000000000000000000000000000";
      s820 <= "0000000000000000000000000000000000";
      s821 <= "0000000000000000000000000000000000";
      s822 <= "0000000000000000000000000000000000";
      s823 <= "0000000000000000000000000000000000";
      s824 <= "0000000000000000000000000000000000";
      s825 <= "0000000000000000000000000000000000";
      s826 <= "0000000000000000000000000000000000";
      s827 <= "0000000000000000000000000000000000";
      s828 <= "0000000000000000000000000000000000";
      s829 <= "0000000000000000000000000000000000";
      s830 <= "0000000000000000000000000000000000";
      s831 <= "0000000000000000000000000000000000";
      s832 <= "0000000000000000000000000000000000";
      s833 <= "0000000000000000000000000000000000";
      s834 <= "0000000000000000000000000000000000";
      s835 <= "0000000000000000000000000000000000";
      s836 <= "0000000000000000000000000000000000";
      s837 <= "0000000000000000000000000000000000";
      s838 <= "0000000000000000000000000000000000";
      s839 <= "0000000000000000000000000000000000";
      s840 <= "0000000000000000000000000000000000";
      s841 <= "0000000000000000000000000000000000";
      s842 <= "0000000000000000000000000000000000";
      s843 <= "0000000000000000000000000000000000";
      s844 <= "0000000000000000000000000000000000";
      s845 <= "0000000000000000000000000000000000";
      s846 <= "0000000000000000000000000000000000";
      s847 <= "0000000000000000000000000000000000";
      s848 <= "0000000000000000000000000000000000";
      s849 <= "0000000000000000000000000000000000";
      s850 <= "0000000000000000000000000000000000";
      s851 <= "0000000000000000000000000000000000";
      s852 <= "0000000000000000000000000000000000";
      s853 <= "0000000000000000000000000000000000";
      s854 <= "0000000000000000000000000000000000";
      s855 <= "0000000000000000000000000000000000";
      s856 <= "0000000000000000000000000000000000";
      s857 <= "0000000000000000000000000000000000";
      s858 <= "0000000000000000000000000000000000";
      s859 <= "0000000000000000000000000000000000";
      s860 <= "0000000000000000000000000000000000";
      s861 <= "0000000000000000000000000000000000";
      s862 <= "0000000000000000000000000000000000";
      s863 <= "0000000000000000000000000000000000";
      s864 <= "0000000000000000000000000000000000";
      s865 <= "0000000000000000000000000000000000";
      s866 <= "0000000000000000000000000000000000";
      s867 <= "0000000000000000000000000000000000";
      s868 <= "0000000000000000000000000000000000";
      s869 <= "0000000000000000000000000000000000";
      s870 <= "0000000000000000000000000000000000";
      s871 <= "0000000000000000000000000000000000";
      s872 <= "0000000000000000000000000000000000";
      s873 <= "0000000000000000000000000000000000";
      s874 <= "0000000000000000000000000000000000";
      s875 <= "0000000000000000000000000000000000";
      s876 <= "0000000000000000000000000000000000";
      s877 <= "0000000000000000000000000000000000";
      s878 <= "0000000000000000000000000000000000";
      s879 <= "0000000000000000000000000000000000";
      s880 <= "0000000000000000000000000000000000";
      s881 <= "0000000000000000000000000000000000";
      s882 <= "0000000000000000000000000000000000";
      s883 <= "0000000000000000000000000000000000";
      s884 <= "0000000000000000000000000000000000";
      s885 <= "0000000000000000000000000000000000";
      s886 <= "0000000000000000000000000000000000";
      s887 <= "0000000000000000000000000000000000";
      s888 <= "0000000000000000000000000000000000";
      s889 <= "0000000000000000000000000000000000";
      s890 <= "0000000000000000000000000000000000";
      s891 <= "0000000000000000000000000000000000";
      s892 <= "0000000000000000000000000000000000";
      s893 <= "0000000000000000000000000000000000";
      s894 <= "0000000000000000000000000000000000";
      s895 <= "0000000000000000000000000000000000";
      s896 <= "0000000000000000000000000000000000";
      s897 <= "0000000000000000000000000000000000";
      s898 <= "0000000000000000000000000000000000";
      s899 <= "0000000000000000000000000000000000";
      s900 <= "0000000000000000000000000000000000";
      s901 <= "0000000000000000000000000000000000";
      s902 <= "0000000000000000000000000000000000";
      s903 <= "0000000000000000000000000000000000";
      s904 <= "0000000000000000000000000000000000";
      s905 <= "0000000000000000000000000000000000";
      s906 <= "0000000000000000000000000000000000";
      s907 <= "0000000000000000000000000000000000";
      s908 <= "0000000000000000000000000000000000";
      s909 <= "0000000000000000000000000000000000";
      s910 <= "0000000000000000000000000000000000";
      s911 <= "0000000000000000000000000000000000";
      s912 <= "0000000000000000000000000000000000";
      s913 <= "0000000000000000000000000000000000";
      s914 <= "0000000000000000000000000000000000";
      s915 <= "0000000000000000000000000000000000";
      s916 <= "0000000000000000000000000000000000";
      s917 <= "0000000000000000000000000000000000";
      s918 <= "0000000000000000000000000000000000";
      s919 <= "0000000000000000000000000000000000";
      s920 <= "0000000000000000000000000000000000";
      s921 <= "0000000000000000000000000000000000";
      s922 <= "0000000000000000000000000000000000";
      s923 <= "0000000000000000000000000000000000";
      s924 <= "0000000000000000000000000000000000";
      s925 <= "0000000000000000000000000000000000";
      s926 <= "0000000000000000000000000000000000";
      s927 <= "0000000000000000000000000000000000";
      s928 <= "0000000000000000000000000000000000";
      s929 <= "0000000000000000000000000000000000";
      s930 <= "0000000000000000000000000000000000";
      s931 <= "0000000000000000000000000000000000";
      s932 <= "0000000000000000000000000000000000";
      s933 <= "0000000000000000000000000000000000";
      s934 <= "0000000000000000000000000000000000";
      s935 <= "0000000000000000000000000000000000";
      s936 <= "0000000000000000000000000000000000";
      s937 <= "0000000000000000000000000000000000";
      s938 <= "0000000000000000000000000000000000";
      s939 <= "0000000000000000000000000000000000";
      s940 <= "0000000000000000000000000000000000";
      s941 <= "0000000000000000000000000000000000";
      s942 <= "0000000000000000000000000000000000";
      s943 <= "0000000000000000000000000000000000";
      s944 <= "0000000000000000000000000000000000";
      s945 <= "0000000000000000000000000000000000";
      s946 <= "0000000000000000000000000000000000";
      s947 <= "0000000000000000000000000000000000";
      s948 <= "0000000000000000000000000000000000";
      s949 <= "0000000000000000000000000000000000";
      s950 <= "0000000000000000000000000000000000";
      s951 <= "0000000000000000000000000000000000";
      s952 <= "0000000000000000000000000000000000";
      s953 <= "0000000000000000000000000000000000";
      s954 <= "0000000000000000000000000000000000";
      s955 <= "0000000000000000000000000000000000";
      s956 <= "0000000000000000000000000000000000";
      s957 <= "0000000000000000000000000000000000";
      s958 <= "0000000000000000000000000000000000";
      s959 <= "0000000000000000000000000000000000";
      s960 <= "0000000000000000000000000000000000";
      s961 <= "0000000000000000000000000000000000";
      s962 <= "0000000000000000000000000000000000";
      s963 <= "0000000000000000000000000000000000";
      s964 <= "0000000000000000000000000000000000";
      s965 <= "0000000000000000000000000000000000";
      s966 <= "0000000000000000000000000000000000";
      s967 <= "0000000000000000000000000000000000";
      s968 <= "0000000000000000000000000000000000";
      s969 <= "0000000000000000000000000000000000";
      s970 <= "0000000000000000000000000000000000";
      s971 <= "0000000000000000000000000000000000";
      s972 <= "0000000000000000000000000000000000";
      s973 <= "0000000000000000000000000000000000";
      s974 <= "0000000000000000000000000000000000";
      s975 <= "0000000000000000000000000000000000";
      s976 <= "0000000000000000000000000000000000";
      s977 <= "0000000000000000000000000000000000";
      s978 <= "0000000000000000000000000000000000";
      s979 <= "0000000000000000000000000000000000";
      s980 <= "0000000000000000000000000000000000";
      s981 <= "0000000000000000000000000000000000";
      s982 <= "0000000000000000000000000000000000";
      s983 <= "0000000000000000000000000000000000";
      s984 <= "0000000000000000000000000000000000";
      s985 <= "0000000000000000000000000000000000";
      s986 <= "0000000000000000000000000000000000";
      s987 <= "0000000000000000000000000000000000";
      s988 <= "0000000000000000000000000000000000";
      s989 <= "0000000000000000000000000000000000";
      s990 <= "0000000000000000000000000000000000";
      s991 <= "0000000000000000000000000000000000";
      s992 <= "0000000000000000000000000000000000";
      s993 <= "0000000000000000000000000000000000";
      s994 <= "0000000000000000000000000000000000";
      s995 <= "0000000000000000000000000000000000";
      s996 <= "0000000000000000000000000000000000";
      s997 <= "0000000000000000000000000000000000";
      s998 <= "0000000000000000000000000000000000";
      s999 <= "0000000000000000000000000000000000";
      s1000 <= "0000000000000000000000000000000000";
      s1001 <= "0000000000000000000000000000000000";
      s1002 <= "0000000000000000000000000000000000";
      s1003 <= "0000000000000000000000000000000000";
      s1004 <= "0000000000000000000000000000000000";
      s1005 <= "0000000000000000000000000000000000";
      s1006 <= "0000000000000000000000000000000000";
      s1007 <= "0000000000000000000000000000000000";
      s1008 <= "0000000000000000000000000000000000";
      s1009 <= "0000000000000000000000000000000000";
      s1010 <= "0000000000000000000000000000000000";
      s1011 <= "0000000000000000000000000000000000";
      s1012 <= "0000000000000000000000000000000000";
      s1013 <= "0000000000000000000000000000000000";
      s1014 <= "0000000000000000000000000000000000";
      s1015 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      s558 <= s557;
      s559 <= s558;
      s560 <= s559;
      s561 <= s560;
      s562 <= s561;
      s563 <= s562;
      s564 <= s563;
      s565 <= s564;
      s566 <= s565;
      s567 <= s566;
      s568 <= s567;
      s569 <= s568;
      s570 <= s569;
      s571 <= s570;
      s572 <= s571;
      s573 <= s572;
      s574 <= s573;
      s575 <= s574;
      s576 <= s575;
      s577 <= s576;
      s578 <= s577;
      s579 <= s578;
      s580 <= s579;
      s581 <= s580;
      s582 <= s581;
      s583 <= s582;
      s584 <= s583;
      s585 <= s584;
      s586 <= s585;
      s587 <= s586;
      s588 <= s587;
      s589 <= s588;
      s590 <= s589;
      s591 <= s590;
      s592 <= s591;
      s593 <= s592;
      s594 <= s593;
      s595 <= s594;
      s596 <= s595;
      s597 <= s596;
      s598 <= s597;
      s599 <= s598;
      s600 <= s599;
      s601 <= s600;
      s602 <= s601;
      s603 <= s602;
      s604 <= s603;
      s605 <= s604;
      s606 <= s605;
      s607 <= s606;
      s608 <= s607;
      s609 <= s608;
      s610 <= s609;
      s611 <= s610;
      s612 <= s611;
      s613 <= s612;
      s614 <= s613;
      s615 <= s614;
      s616 <= s615;
      s617 <= s616;
      s618 <= s617;
      s619 <= s618;
      s620 <= s619;
      s621 <= s620;
      s622 <= s621;
      s623 <= s622;
      s624 <= s623;
      s625 <= s624;
      s626 <= s625;
      s627 <= s626;
      s628 <= s627;
      s629 <= s628;
      s630 <= s629;
      s631 <= s630;
      s632 <= s631;
      s633 <= s632;
      s634 <= s633;
      s635 <= s634;
      s636 <= s635;
      s637 <= s636;
      s638 <= s637;
      s639 <= s638;
      s640 <= s639;
      s641 <= s640;
      s642 <= s641;
      s643 <= s642;
      s644 <= s643;
      s645 <= s644;
      s646 <= s645;
      s647 <= s646;
      s648 <= s647;
      s649 <= s648;
      s650 <= s649;
      s651 <= s650;
      s652 <= s651;
      s653 <= s652;
      s654 <= s653;
      s655 <= s654;
      s656 <= s655;
      s657 <= s656;
      s658 <= s657;
      s659 <= s658;
      s660 <= s659;
      s661 <= s660;
      s662 <= s661;
      s663 <= s662;
      s664 <= s663;
      s665 <= s664;
      s666 <= s665;
      s667 <= s666;
      s668 <= s667;
      s669 <= s668;
      s670 <= s669;
      s671 <= s670;
      s672 <= s671;
      s673 <= s672;
      s674 <= s673;
      s675 <= s674;
      s676 <= s675;
      s677 <= s676;
      s678 <= s677;
      s679 <= s678;
      s680 <= s679;
      s681 <= s680;
      s682 <= s681;
      s683 <= s682;
      s684 <= s683;
      s685 <= s684;
      s686 <= s685;
      s687 <= s686;
      s688 <= s687;
      s689 <= s688;
      s690 <= s689;
      s691 <= s690;
      s692 <= s691;
      s693 <= s692;
      s694 <= s693;
      s695 <= s694;
      s696 <= s695;
      s697 <= s696;
      s698 <= s697;
      s699 <= s698;
      s700 <= s699;
      s701 <= s700;
      s702 <= s701;
      s703 <= s702;
      s704 <= s703;
      s705 <= s704;
      s706 <= s705;
      s707 <= s706;
      s708 <= s707;
      s709 <= s708;
      s710 <= s709;
      s711 <= s710;
      s712 <= s711;
      s713 <= s712;
      s714 <= s713;
      s715 <= s714;
      s716 <= s715;
      s717 <= s716;
      s718 <= s717;
      s719 <= s718;
      s720 <= s719;
      s721 <= s720;
      s722 <= s721;
      s723 <= s722;
      s724 <= s723;
      s725 <= s724;
      s726 <= s725;
      s727 <= s726;
      s728 <= s727;
      s729 <= s728;
      s730 <= s729;
      s731 <= s730;
      s732 <= s731;
      s733 <= s732;
      s734 <= s733;
      s735 <= s734;
      s736 <= s735;
      s737 <= s736;
      s738 <= s737;
      s739 <= s738;
      s740 <= s739;
      s741 <= s740;
      s742 <= s741;
      s743 <= s742;
      s744 <= s743;
      s745 <= s744;
      s746 <= s745;
      s747 <= s746;
      s748 <= s747;
      s749 <= s748;
      s750 <= s749;
      s751 <= s750;
      s752 <= s751;
      s753 <= s752;
      s754 <= s753;
      s755 <= s754;
      s756 <= s755;
      s757 <= s756;
      s758 <= s757;
      s759 <= s758;
      s760 <= s759;
      s761 <= s760;
      s762 <= s761;
      s763 <= s762;
      s764 <= s763;
      s765 <= s764;
      s766 <= s765;
      s767 <= s766;
      s768 <= s767;
      s769 <= s768;
      s770 <= s769;
      s771 <= s770;
      s772 <= s771;
      s773 <= s772;
      s774 <= s773;
      s775 <= s774;
      s776 <= s775;
      s777 <= s776;
      s778 <= s777;
      s779 <= s778;
      s780 <= s779;
      s781 <= s780;
      s782 <= s781;
      s783 <= s782;
      s784 <= s783;
      s785 <= s784;
      s786 <= s785;
      s787 <= s786;
      s788 <= s787;
      s789 <= s788;
      s790 <= s789;
      s791 <= s790;
      s792 <= s791;
      s793 <= s792;
      s794 <= s793;
      s795 <= s794;
      s796 <= s795;
      s797 <= s796;
      s798 <= s797;
      s799 <= s798;
      s800 <= s799;
      s801 <= s800;
      s802 <= s801;
      s803 <= s802;
      s804 <= s803;
      s805 <= s804;
      s806 <= s805;
      s807 <= s806;
      s808 <= s807;
      s809 <= s808;
      s810 <= s809;
      s811 <= s810;
      s812 <= s811;
      s813 <= s812;
      s814 <= s813;
      s815 <= s814;
      s816 <= s815;
      s817 <= s816;
      s818 <= s817;
      s819 <= s818;
      s820 <= s819;
      s821 <= s820;
      s822 <= s821;
      s823 <= s822;
      s824 <= s823;
      s825 <= s824;
      s826 <= s825;
      s827 <= s826;
      s828 <= s827;
      s829 <= s828;
      s830 <= s829;
      s831 <= s830;
      s832 <= s831;
      s833 <= s832;
      s834 <= s833;
      s835 <= s834;
      s836 <= s835;
      s837 <= s836;
      s838 <= s837;
      s839 <= s838;
      s840 <= s839;
      s841 <= s840;
      s842 <= s841;
      s843 <= s842;
      s844 <= s843;
      s845 <= s844;
      s846 <= s845;
      s847 <= s846;
      s848 <= s847;
      s849 <= s848;
      s850 <= s849;
      s851 <= s850;
      s852 <= s851;
      s853 <= s852;
      s854 <= s853;
      s855 <= s854;
      s856 <= s855;
      s857 <= s856;
      s858 <= s857;
      s859 <= s858;
      s860 <= s859;
      s861 <= s860;
      s862 <= s861;
      s863 <= s862;
      s864 <= s863;
      s865 <= s864;
      s866 <= s865;
      s867 <= s866;
      s868 <= s867;
      s869 <= s868;
      s870 <= s869;
      s871 <= s870;
      s872 <= s871;
      s873 <= s872;
      s874 <= s873;
      s875 <= s874;
      s876 <= s875;
      s877 <= s876;
      s878 <= s877;
      s879 <= s878;
      s880 <= s879;
      s881 <= s880;
      s882 <= s881;
      s883 <= s882;
      s884 <= s883;
      s885 <= s884;
      s886 <= s885;
      s887 <= s886;
      s888 <= s887;
      s889 <= s888;
      s890 <= s889;
      s891 <= s890;
      s892 <= s891;
      s893 <= s892;
      s894 <= s893;
      s895 <= s894;
      s896 <= s895;
      s897 <= s896;
      s898 <= s897;
      s899 <= s898;
      s900 <= s899;
      s901 <= s900;
      s902 <= s901;
      s903 <= s902;
      s904 <= s903;
      s905 <= s904;
      s906 <= s905;
      s907 <= s906;
      s908 <= s907;
      s909 <= s908;
      s910 <= s909;
      s911 <= s910;
      s912 <= s911;
      s913 <= s912;
      s914 <= s913;
      s915 <= s914;
      s916 <= s915;
      s917 <= s916;
      s918 <= s917;
      s919 <= s918;
      s920 <= s919;
      s921 <= s920;
      s922 <= s921;
      s923 <= s922;
      s924 <= s923;
      s925 <= s924;
      s926 <= s925;
      s927 <= s926;
      s928 <= s927;
      s929 <= s928;
      s930 <= s929;
      s931 <= s930;
      s932 <= s931;
      s933 <= s932;
      s934 <= s933;
      s935 <= s934;
      s936 <= s935;
      s937 <= s936;
      s938 <= s937;
      s939 <= s938;
      s940 <= s939;
      s941 <= s940;
      s942 <= s941;
      s943 <= s942;
      s944 <= s943;
      s945 <= s944;
      s946 <= s945;
      s947 <= s946;
      s948 <= s947;
      s949 <= s948;
      s950 <= s949;
      s951 <= s950;
      s952 <= s951;
      s953 <= s952;
      s954 <= s953;
      s955 <= s954;
      s956 <= s955;
      s957 <= s956;
      s958 <= s957;
      s959 <= s958;
      s960 <= s959;
      s961 <= s960;
      s962 <= s961;
      s963 <= s962;
      s964 <= s963;
      s965 <= s964;
      s966 <= s965;
      s967 <= s966;
      s968 <= s967;
      s969 <= s968;
      s970 <= s969;
      s971 <= s970;
      s972 <= s971;
      s973 <= s972;
      s974 <= s973;
      s975 <= s974;
      s976 <= s975;
      s977 <= s976;
      s978 <= s977;
      s979 <= s978;
      s980 <= s979;
      s981 <= s980;
      s982 <= s981;
      s983 <= s982;
      s984 <= s983;
      s985 <= s984;
      s986 <= s985;
      s987 <= s986;
      s988 <= s987;
      s989 <= s988;
      s990 <= s989;
      s991 <= s990;
      s992 <= s991;
      s993 <= s992;
      s994 <= s993;
      s995 <= s994;
      s996 <= s995;
      s997 <= s996;
      s998 <= s997;
      s999 <= s998;
      s1000 <= s999;
      s1001 <= s1000;
      s1002 <= s1001;
      s1003 <= s1002;
      s1004 <= s1003;
      s1005 <= s1004;
      s1006 <= s1005;
      s1007 <= s1006;
      s1008 <= s1007;
      s1009 <= s1008;
      s1010 <= s1009;
      s1011 <= s1010;
      s1012 <= s1011;
      s1013 <= s1012;
      s1014 <= s1013;
      s1015 <= s1014;
      Y <= s1015;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1081_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1081 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1081_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1081_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
signal s558 : std_logic_vector(33 downto 0) := (others => '0');
signal s559 : std_logic_vector(33 downto 0) := (others => '0');
signal s560 : std_logic_vector(33 downto 0) := (others => '0');
signal s561 : std_logic_vector(33 downto 0) := (others => '0');
signal s562 : std_logic_vector(33 downto 0) := (others => '0');
signal s563 : std_logic_vector(33 downto 0) := (others => '0');
signal s564 : std_logic_vector(33 downto 0) := (others => '0');
signal s565 : std_logic_vector(33 downto 0) := (others => '0');
signal s566 : std_logic_vector(33 downto 0) := (others => '0');
signal s567 : std_logic_vector(33 downto 0) := (others => '0');
signal s568 : std_logic_vector(33 downto 0) := (others => '0');
signal s569 : std_logic_vector(33 downto 0) := (others => '0');
signal s570 : std_logic_vector(33 downto 0) := (others => '0');
signal s571 : std_logic_vector(33 downto 0) := (others => '0');
signal s572 : std_logic_vector(33 downto 0) := (others => '0');
signal s573 : std_logic_vector(33 downto 0) := (others => '0');
signal s574 : std_logic_vector(33 downto 0) := (others => '0');
signal s575 : std_logic_vector(33 downto 0) := (others => '0');
signal s576 : std_logic_vector(33 downto 0) := (others => '0');
signal s577 : std_logic_vector(33 downto 0) := (others => '0');
signal s578 : std_logic_vector(33 downto 0) := (others => '0');
signal s579 : std_logic_vector(33 downto 0) := (others => '0');
signal s580 : std_logic_vector(33 downto 0) := (others => '0');
signal s581 : std_logic_vector(33 downto 0) := (others => '0');
signal s582 : std_logic_vector(33 downto 0) := (others => '0');
signal s583 : std_logic_vector(33 downto 0) := (others => '0');
signal s584 : std_logic_vector(33 downto 0) := (others => '0');
signal s585 : std_logic_vector(33 downto 0) := (others => '0');
signal s586 : std_logic_vector(33 downto 0) := (others => '0');
signal s587 : std_logic_vector(33 downto 0) := (others => '0');
signal s588 : std_logic_vector(33 downto 0) := (others => '0');
signal s589 : std_logic_vector(33 downto 0) := (others => '0');
signal s590 : std_logic_vector(33 downto 0) := (others => '0');
signal s591 : std_logic_vector(33 downto 0) := (others => '0');
signal s592 : std_logic_vector(33 downto 0) := (others => '0');
signal s593 : std_logic_vector(33 downto 0) := (others => '0');
signal s594 : std_logic_vector(33 downto 0) := (others => '0');
signal s595 : std_logic_vector(33 downto 0) := (others => '0');
signal s596 : std_logic_vector(33 downto 0) := (others => '0');
signal s597 : std_logic_vector(33 downto 0) := (others => '0');
signal s598 : std_logic_vector(33 downto 0) := (others => '0');
signal s599 : std_logic_vector(33 downto 0) := (others => '0');
signal s600 : std_logic_vector(33 downto 0) := (others => '0');
signal s601 : std_logic_vector(33 downto 0) := (others => '0');
signal s602 : std_logic_vector(33 downto 0) := (others => '0');
signal s603 : std_logic_vector(33 downto 0) := (others => '0');
signal s604 : std_logic_vector(33 downto 0) := (others => '0');
signal s605 : std_logic_vector(33 downto 0) := (others => '0');
signal s606 : std_logic_vector(33 downto 0) := (others => '0');
signal s607 : std_logic_vector(33 downto 0) := (others => '0');
signal s608 : std_logic_vector(33 downto 0) := (others => '0');
signal s609 : std_logic_vector(33 downto 0) := (others => '0');
signal s610 : std_logic_vector(33 downto 0) := (others => '0');
signal s611 : std_logic_vector(33 downto 0) := (others => '0');
signal s612 : std_logic_vector(33 downto 0) := (others => '0');
signal s613 : std_logic_vector(33 downto 0) := (others => '0');
signal s614 : std_logic_vector(33 downto 0) := (others => '0');
signal s615 : std_logic_vector(33 downto 0) := (others => '0');
signal s616 : std_logic_vector(33 downto 0) := (others => '0');
signal s617 : std_logic_vector(33 downto 0) := (others => '0');
signal s618 : std_logic_vector(33 downto 0) := (others => '0');
signal s619 : std_logic_vector(33 downto 0) := (others => '0');
signal s620 : std_logic_vector(33 downto 0) := (others => '0');
signal s621 : std_logic_vector(33 downto 0) := (others => '0');
signal s622 : std_logic_vector(33 downto 0) := (others => '0');
signal s623 : std_logic_vector(33 downto 0) := (others => '0');
signal s624 : std_logic_vector(33 downto 0) := (others => '0');
signal s625 : std_logic_vector(33 downto 0) := (others => '0');
signal s626 : std_logic_vector(33 downto 0) := (others => '0');
signal s627 : std_logic_vector(33 downto 0) := (others => '0');
signal s628 : std_logic_vector(33 downto 0) := (others => '0');
signal s629 : std_logic_vector(33 downto 0) := (others => '0');
signal s630 : std_logic_vector(33 downto 0) := (others => '0');
signal s631 : std_logic_vector(33 downto 0) := (others => '0');
signal s632 : std_logic_vector(33 downto 0) := (others => '0');
signal s633 : std_logic_vector(33 downto 0) := (others => '0');
signal s634 : std_logic_vector(33 downto 0) := (others => '0');
signal s635 : std_logic_vector(33 downto 0) := (others => '0');
signal s636 : std_logic_vector(33 downto 0) := (others => '0');
signal s637 : std_logic_vector(33 downto 0) := (others => '0');
signal s638 : std_logic_vector(33 downto 0) := (others => '0');
signal s639 : std_logic_vector(33 downto 0) := (others => '0');
signal s640 : std_logic_vector(33 downto 0) := (others => '0');
signal s641 : std_logic_vector(33 downto 0) := (others => '0');
signal s642 : std_logic_vector(33 downto 0) := (others => '0');
signal s643 : std_logic_vector(33 downto 0) := (others => '0');
signal s644 : std_logic_vector(33 downto 0) := (others => '0');
signal s645 : std_logic_vector(33 downto 0) := (others => '0');
signal s646 : std_logic_vector(33 downto 0) := (others => '0');
signal s647 : std_logic_vector(33 downto 0) := (others => '0');
signal s648 : std_logic_vector(33 downto 0) := (others => '0');
signal s649 : std_logic_vector(33 downto 0) := (others => '0');
signal s650 : std_logic_vector(33 downto 0) := (others => '0');
signal s651 : std_logic_vector(33 downto 0) := (others => '0');
signal s652 : std_logic_vector(33 downto 0) := (others => '0');
signal s653 : std_logic_vector(33 downto 0) := (others => '0');
signal s654 : std_logic_vector(33 downto 0) := (others => '0');
signal s655 : std_logic_vector(33 downto 0) := (others => '0');
signal s656 : std_logic_vector(33 downto 0) := (others => '0');
signal s657 : std_logic_vector(33 downto 0) := (others => '0');
signal s658 : std_logic_vector(33 downto 0) := (others => '0');
signal s659 : std_logic_vector(33 downto 0) := (others => '0');
signal s660 : std_logic_vector(33 downto 0) := (others => '0');
signal s661 : std_logic_vector(33 downto 0) := (others => '0');
signal s662 : std_logic_vector(33 downto 0) := (others => '0');
signal s663 : std_logic_vector(33 downto 0) := (others => '0');
signal s664 : std_logic_vector(33 downto 0) := (others => '0');
signal s665 : std_logic_vector(33 downto 0) := (others => '0');
signal s666 : std_logic_vector(33 downto 0) := (others => '0');
signal s667 : std_logic_vector(33 downto 0) := (others => '0');
signal s668 : std_logic_vector(33 downto 0) := (others => '0');
signal s669 : std_logic_vector(33 downto 0) := (others => '0');
signal s670 : std_logic_vector(33 downto 0) := (others => '0');
signal s671 : std_logic_vector(33 downto 0) := (others => '0');
signal s672 : std_logic_vector(33 downto 0) := (others => '0');
signal s673 : std_logic_vector(33 downto 0) := (others => '0');
signal s674 : std_logic_vector(33 downto 0) := (others => '0');
signal s675 : std_logic_vector(33 downto 0) := (others => '0');
signal s676 : std_logic_vector(33 downto 0) := (others => '0');
signal s677 : std_logic_vector(33 downto 0) := (others => '0');
signal s678 : std_logic_vector(33 downto 0) := (others => '0');
signal s679 : std_logic_vector(33 downto 0) := (others => '0');
signal s680 : std_logic_vector(33 downto 0) := (others => '0');
signal s681 : std_logic_vector(33 downto 0) := (others => '0');
signal s682 : std_logic_vector(33 downto 0) := (others => '0');
signal s683 : std_logic_vector(33 downto 0) := (others => '0');
signal s684 : std_logic_vector(33 downto 0) := (others => '0');
signal s685 : std_logic_vector(33 downto 0) := (others => '0');
signal s686 : std_logic_vector(33 downto 0) := (others => '0');
signal s687 : std_logic_vector(33 downto 0) := (others => '0');
signal s688 : std_logic_vector(33 downto 0) := (others => '0');
signal s689 : std_logic_vector(33 downto 0) := (others => '0');
signal s690 : std_logic_vector(33 downto 0) := (others => '0');
signal s691 : std_logic_vector(33 downto 0) := (others => '0');
signal s692 : std_logic_vector(33 downto 0) := (others => '0');
signal s693 : std_logic_vector(33 downto 0) := (others => '0');
signal s694 : std_logic_vector(33 downto 0) := (others => '0');
signal s695 : std_logic_vector(33 downto 0) := (others => '0');
signal s696 : std_logic_vector(33 downto 0) := (others => '0');
signal s697 : std_logic_vector(33 downto 0) := (others => '0');
signal s698 : std_logic_vector(33 downto 0) := (others => '0');
signal s699 : std_logic_vector(33 downto 0) := (others => '0');
signal s700 : std_logic_vector(33 downto 0) := (others => '0');
signal s701 : std_logic_vector(33 downto 0) := (others => '0');
signal s702 : std_logic_vector(33 downto 0) := (others => '0');
signal s703 : std_logic_vector(33 downto 0) := (others => '0');
signal s704 : std_logic_vector(33 downto 0) := (others => '0');
signal s705 : std_logic_vector(33 downto 0) := (others => '0');
signal s706 : std_logic_vector(33 downto 0) := (others => '0');
signal s707 : std_logic_vector(33 downto 0) := (others => '0');
signal s708 : std_logic_vector(33 downto 0) := (others => '0');
signal s709 : std_logic_vector(33 downto 0) := (others => '0');
signal s710 : std_logic_vector(33 downto 0) := (others => '0');
signal s711 : std_logic_vector(33 downto 0) := (others => '0');
signal s712 : std_logic_vector(33 downto 0) := (others => '0');
signal s713 : std_logic_vector(33 downto 0) := (others => '0');
signal s714 : std_logic_vector(33 downto 0) := (others => '0');
signal s715 : std_logic_vector(33 downto 0) := (others => '0');
signal s716 : std_logic_vector(33 downto 0) := (others => '0');
signal s717 : std_logic_vector(33 downto 0) := (others => '0');
signal s718 : std_logic_vector(33 downto 0) := (others => '0');
signal s719 : std_logic_vector(33 downto 0) := (others => '0');
signal s720 : std_logic_vector(33 downto 0) := (others => '0');
signal s721 : std_logic_vector(33 downto 0) := (others => '0');
signal s722 : std_logic_vector(33 downto 0) := (others => '0');
signal s723 : std_logic_vector(33 downto 0) := (others => '0');
signal s724 : std_logic_vector(33 downto 0) := (others => '0');
signal s725 : std_logic_vector(33 downto 0) := (others => '0');
signal s726 : std_logic_vector(33 downto 0) := (others => '0');
signal s727 : std_logic_vector(33 downto 0) := (others => '0');
signal s728 : std_logic_vector(33 downto 0) := (others => '0');
signal s729 : std_logic_vector(33 downto 0) := (others => '0');
signal s730 : std_logic_vector(33 downto 0) := (others => '0');
signal s731 : std_logic_vector(33 downto 0) := (others => '0');
signal s732 : std_logic_vector(33 downto 0) := (others => '0');
signal s733 : std_logic_vector(33 downto 0) := (others => '0');
signal s734 : std_logic_vector(33 downto 0) := (others => '0');
signal s735 : std_logic_vector(33 downto 0) := (others => '0');
signal s736 : std_logic_vector(33 downto 0) := (others => '0');
signal s737 : std_logic_vector(33 downto 0) := (others => '0');
signal s738 : std_logic_vector(33 downto 0) := (others => '0');
signal s739 : std_logic_vector(33 downto 0) := (others => '0');
signal s740 : std_logic_vector(33 downto 0) := (others => '0');
signal s741 : std_logic_vector(33 downto 0) := (others => '0');
signal s742 : std_logic_vector(33 downto 0) := (others => '0');
signal s743 : std_logic_vector(33 downto 0) := (others => '0');
signal s744 : std_logic_vector(33 downto 0) := (others => '0');
signal s745 : std_logic_vector(33 downto 0) := (others => '0');
signal s746 : std_logic_vector(33 downto 0) := (others => '0');
signal s747 : std_logic_vector(33 downto 0) := (others => '0');
signal s748 : std_logic_vector(33 downto 0) := (others => '0');
signal s749 : std_logic_vector(33 downto 0) := (others => '0');
signal s750 : std_logic_vector(33 downto 0) := (others => '0');
signal s751 : std_logic_vector(33 downto 0) := (others => '0');
signal s752 : std_logic_vector(33 downto 0) := (others => '0');
signal s753 : std_logic_vector(33 downto 0) := (others => '0');
signal s754 : std_logic_vector(33 downto 0) := (others => '0');
signal s755 : std_logic_vector(33 downto 0) := (others => '0');
signal s756 : std_logic_vector(33 downto 0) := (others => '0');
signal s757 : std_logic_vector(33 downto 0) := (others => '0');
signal s758 : std_logic_vector(33 downto 0) := (others => '0');
signal s759 : std_logic_vector(33 downto 0) := (others => '0');
signal s760 : std_logic_vector(33 downto 0) := (others => '0');
signal s761 : std_logic_vector(33 downto 0) := (others => '0');
signal s762 : std_logic_vector(33 downto 0) := (others => '0');
signal s763 : std_logic_vector(33 downto 0) := (others => '0');
signal s764 : std_logic_vector(33 downto 0) := (others => '0');
signal s765 : std_logic_vector(33 downto 0) := (others => '0');
signal s766 : std_logic_vector(33 downto 0) := (others => '0');
signal s767 : std_logic_vector(33 downto 0) := (others => '0');
signal s768 : std_logic_vector(33 downto 0) := (others => '0');
signal s769 : std_logic_vector(33 downto 0) := (others => '0');
signal s770 : std_logic_vector(33 downto 0) := (others => '0');
signal s771 : std_logic_vector(33 downto 0) := (others => '0');
signal s772 : std_logic_vector(33 downto 0) := (others => '0');
signal s773 : std_logic_vector(33 downto 0) := (others => '0');
signal s774 : std_logic_vector(33 downto 0) := (others => '0');
signal s775 : std_logic_vector(33 downto 0) := (others => '0');
signal s776 : std_logic_vector(33 downto 0) := (others => '0');
signal s777 : std_logic_vector(33 downto 0) := (others => '0');
signal s778 : std_logic_vector(33 downto 0) := (others => '0');
signal s779 : std_logic_vector(33 downto 0) := (others => '0');
signal s780 : std_logic_vector(33 downto 0) := (others => '0');
signal s781 : std_logic_vector(33 downto 0) := (others => '0');
signal s782 : std_logic_vector(33 downto 0) := (others => '0');
signal s783 : std_logic_vector(33 downto 0) := (others => '0');
signal s784 : std_logic_vector(33 downto 0) := (others => '0');
signal s785 : std_logic_vector(33 downto 0) := (others => '0');
signal s786 : std_logic_vector(33 downto 0) := (others => '0');
signal s787 : std_logic_vector(33 downto 0) := (others => '0');
signal s788 : std_logic_vector(33 downto 0) := (others => '0');
signal s789 : std_logic_vector(33 downto 0) := (others => '0');
signal s790 : std_logic_vector(33 downto 0) := (others => '0');
signal s791 : std_logic_vector(33 downto 0) := (others => '0');
signal s792 : std_logic_vector(33 downto 0) := (others => '0');
signal s793 : std_logic_vector(33 downto 0) := (others => '0');
signal s794 : std_logic_vector(33 downto 0) := (others => '0');
signal s795 : std_logic_vector(33 downto 0) := (others => '0');
signal s796 : std_logic_vector(33 downto 0) := (others => '0');
signal s797 : std_logic_vector(33 downto 0) := (others => '0');
signal s798 : std_logic_vector(33 downto 0) := (others => '0');
signal s799 : std_logic_vector(33 downto 0) := (others => '0');
signal s800 : std_logic_vector(33 downto 0) := (others => '0');
signal s801 : std_logic_vector(33 downto 0) := (others => '0');
signal s802 : std_logic_vector(33 downto 0) := (others => '0');
signal s803 : std_logic_vector(33 downto 0) := (others => '0');
signal s804 : std_logic_vector(33 downto 0) := (others => '0');
signal s805 : std_logic_vector(33 downto 0) := (others => '0');
signal s806 : std_logic_vector(33 downto 0) := (others => '0');
signal s807 : std_logic_vector(33 downto 0) := (others => '0');
signal s808 : std_logic_vector(33 downto 0) := (others => '0');
signal s809 : std_logic_vector(33 downto 0) := (others => '0');
signal s810 : std_logic_vector(33 downto 0) := (others => '0');
signal s811 : std_logic_vector(33 downto 0) := (others => '0');
signal s812 : std_logic_vector(33 downto 0) := (others => '0');
signal s813 : std_logic_vector(33 downto 0) := (others => '0');
signal s814 : std_logic_vector(33 downto 0) := (others => '0');
signal s815 : std_logic_vector(33 downto 0) := (others => '0');
signal s816 : std_logic_vector(33 downto 0) := (others => '0');
signal s817 : std_logic_vector(33 downto 0) := (others => '0');
signal s818 : std_logic_vector(33 downto 0) := (others => '0');
signal s819 : std_logic_vector(33 downto 0) := (others => '0');
signal s820 : std_logic_vector(33 downto 0) := (others => '0');
signal s821 : std_logic_vector(33 downto 0) := (others => '0');
signal s822 : std_logic_vector(33 downto 0) := (others => '0');
signal s823 : std_logic_vector(33 downto 0) := (others => '0');
signal s824 : std_logic_vector(33 downto 0) := (others => '0');
signal s825 : std_logic_vector(33 downto 0) := (others => '0');
signal s826 : std_logic_vector(33 downto 0) := (others => '0');
signal s827 : std_logic_vector(33 downto 0) := (others => '0');
signal s828 : std_logic_vector(33 downto 0) := (others => '0');
signal s829 : std_logic_vector(33 downto 0) := (others => '0');
signal s830 : std_logic_vector(33 downto 0) := (others => '0');
signal s831 : std_logic_vector(33 downto 0) := (others => '0');
signal s832 : std_logic_vector(33 downto 0) := (others => '0');
signal s833 : std_logic_vector(33 downto 0) := (others => '0');
signal s834 : std_logic_vector(33 downto 0) := (others => '0');
signal s835 : std_logic_vector(33 downto 0) := (others => '0');
signal s836 : std_logic_vector(33 downto 0) := (others => '0');
signal s837 : std_logic_vector(33 downto 0) := (others => '0');
signal s838 : std_logic_vector(33 downto 0) := (others => '0');
signal s839 : std_logic_vector(33 downto 0) := (others => '0');
signal s840 : std_logic_vector(33 downto 0) := (others => '0');
signal s841 : std_logic_vector(33 downto 0) := (others => '0');
signal s842 : std_logic_vector(33 downto 0) := (others => '0');
signal s843 : std_logic_vector(33 downto 0) := (others => '0');
signal s844 : std_logic_vector(33 downto 0) := (others => '0');
signal s845 : std_logic_vector(33 downto 0) := (others => '0');
signal s846 : std_logic_vector(33 downto 0) := (others => '0');
signal s847 : std_logic_vector(33 downto 0) := (others => '0');
signal s848 : std_logic_vector(33 downto 0) := (others => '0');
signal s849 : std_logic_vector(33 downto 0) := (others => '0');
signal s850 : std_logic_vector(33 downto 0) := (others => '0');
signal s851 : std_logic_vector(33 downto 0) := (others => '0');
signal s852 : std_logic_vector(33 downto 0) := (others => '0');
signal s853 : std_logic_vector(33 downto 0) := (others => '0');
signal s854 : std_logic_vector(33 downto 0) := (others => '0');
signal s855 : std_logic_vector(33 downto 0) := (others => '0');
signal s856 : std_logic_vector(33 downto 0) := (others => '0');
signal s857 : std_logic_vector(33 downto 0) := (others => '0');
signal s858 : std_logic_vector(33 downto 0) := (others => '0');
signal s859 : std_logic_vector(33 downto 0) := (others => '0');
signal s860 : std_logic_vector(33 downto 0) := (others => '0');
signal s861 : std_logic_vector(33 downto 0) := (others => '0');
signal s862 : std_logic_vector(33 downto 0) := (others => '0');
signal s863 : std_logic_vector(33 downto 0) := (others => '0');
signal s864 : std_logic_vector(33 downto 0) := (others => '0');
signal s865 : std_logic_vector(33 downto 0) := (others => '0');
signal s866 : std_logic_vector(33 downto 0) := (others => '0');
signal s867 : std_logic_vector(33 downto 0) := (others => '0');
signal s868 : std_logic_vector(33 downto 0) := (others => '0');
signal s869 : std_logic_vector(33 downto 0) := (others => '0');
signal s870 : std_logic_vector(33 downto 0) := (others => '0');
signal s871 : std_logic_vector(33 downto 0) := (others => '0');
signal s872 : std_logic_vector(33 downto 0) := (others => '0');
signal s873 : std_logic_vector(33 downto 0) := (others => '0');
signal s874 : std_logic_vector(33 downto 0) := (others => '0');
signal s875 : std_logic_vector(33 downto 0) := (others => '0');
signal s876 : std_logic_vector(33 downto 0) := (others => '0');
signal s877 : std_logic_vector(33 downto 0) := (others => '0');
signal s878 : std_logic_vector(33 downto 0) := (others => '0');
signal s879 : std_logic_vector(33 downto 0) := (others => '0');
signal s880 : std_logic_vector(33 downto 0) := (others => '0');
signal s881 : std_logic_vector(33 downto 0) := (others => '0');
signal s882 : std_logic_vector(33 downto 0) := (others => '0');
signal s883 : std_logic_vector(33 downto 0) := (others => '0');
signal s884 : std_logic_vector(33 downto 0) := (others => '0');
signal s885 : std_logic_vector(33 downto 0) := (others => '0');
signal s886 : std_logic_vector(33 downto 0) := (others => '0');
signal s887 : std_logic_vector(33 downto 0) := (others => '0');
signal s888 : std_logic_vector(33 downto 0) := (others => '0');
signal s889 : std_logic_vector(33 downto 0) := (others => '0');
signal s890 : std_logic_vector(33 downto 0) := (others => '0');
signal s891 : std_logic_vector(33 downto 0) := (others => '0');
signal s892 : std_logic_vector(33 downto 0) := (others => '0');
signal s893 : std_logic_vector(33 downto 0) := (others => '0');
signal s894 : std_logic_vector(33 downto 0) := (others => '0');
signal s895 : std_logic_vector(33 downto 0) := (others => '0');
signal s896 : std_logic_vector(33 downto 0) := (others => '0');
signal s897 : std_logic_vector(33 downto 0) := (others => '0');
signal s898 : std_logic_vector(33 downto 0) := (others => '0');
signal s899 : std_logic_vector(33 downto 0) := (others => '0');
signal s900 : std_logic_vector(33 downto 0) := (others => '0');
signal s901 : std_logic_vector(33 downto 0) := (others => '0');
signal s902 : std_logic_vector(33 downto 0) := (others => '0');
signal s903 : std_logic_vector(33 downto 0) := (others => '0');
signal s904 : std_logic_vector(33 downto 0) := (others => '0');
signal s905 : std_logic_vector(33 downto 0) := (others => '0');
signal s906 : std_logic_vector(33 downto 0) := (others => '0');
signal s907 : std_logic_vector(33 downto 0) := (others => '0');
signal s908 : std_logic_vector(33 downto 0) := (others => '0');
signal s909 : std_logic_vector(33 downto 0) := (others => '0');
signal s910 : std_logic_vector(33 downto 0) := (others => '0');
signal s911 : std_logic_vector(33 downto 0) := (others => '0');
signal s912 : std_logic_vector(33 downto 0) := (others => '0');
signal s913 : std_logic_vector(33 downto 0) := (others => '0');
signal s914 : std_logic_vector(33 downto 0) := (others => '0');
signal s915 : std_logic_vector(33 downto 0) := (others => '0');
signal s916 : std_logic_vector(33 downto 0) := (others => '0');
signal s917 : std_logic_vector(33 downto 0) := (others => '0');
signal s918 : std_logic_vector(33 downto 0) := (others => '0');
signal s919 : std_logic_vector(33 downto 0) := (others => '0');
signal s920 : std_logic_vector(33 downto 0) := (others => '0');
signal s921 : std_logic_vector(33 downto 0) := (others => '0');
signal s922 : std_logic_vector(33 downto 0) := (others => '0');
signal s923 : std_logic_vector(33 downto 0) := (others => '0');
signal s924 : std_logic_vector(33 downto 0) := (others => '0');
signal s925 : std_logic_vector(33 downto 0) := (others => '0');
signal s926 : std_logic_vector(33 downto 0) := (others => '0');
signal s927 : std_logic_vector(33 downto 0) := (others => '0');
signal s928 : std_logic_vector(33 downto 0) := (others => '0');
signal s929 : std_logic_vector(33 downto 0) := (others => '0');
signal s930 : std_logic_vector(33 downto 0) := (others => '0');
signal s931 : std_logic_vector(33 downto 0) := (others => '0');
signal s932 : std_logic_vector(33 downto 0) := (others => '0');
signal s933 : std_logic_vector(33 downto 0) := (others => '0');
signal s934 : std_logic_vector(33 downto 0) := (others => '0');
signal s935 : std_logic_vector(33 downto 0) := (others => '0');
signal s936 : std_logic_vector(33 downto 0) := (others => '0');
signal s937 : std_logic_vector(33 downto 0) := (others => '0');
signal s938 : std_logic_vector(33 downto 0) := (others => '0');
signal s939 : std_logic_vector(33 downto 0) := (others => '0');
signal s940 : std_logic_vector(33 downto 0) := (others => '0');
signal s941 : std_logic_vector(33 downto 0) := (others => '0');
signal s942 : std_logic_vector(33 downto 0) := (others => '0');
signal s943 : std_logic_vector(33 downto 0) := (others => '0');
signal s944 : std_logic_vector(33 downto 0) := (others => '0');
signal s945 : std_logic_vector(33 downto 0) := (others => '0');
signal s946 : std_logic_vector(33 downto 0) := (others => '0');
signal s947 : std_logic_vector(33 downto 0) := (others => '0');
signal s948 : std_logic_vector(33 downto 0) := (others => '0');
signal s949 : std_logic_vector(33 downto 0) := (others => '0');
signal s950 : std_logic_vector(33 downto 0) := (others => '0');
signal s951 : std_logic_vector(33 downto 0) := (others => '0');
signal s952 : std_logic_vector(33 downto 0) := (others => '0');
signal s953 : std_logic_vector(33 downto 0) := (others => '0');
signal s954 : std_logic_vector(33 downto 0) := (others => '0');
signal s955 : std_logic_vector(33 downto 0) := (others => '0');
signal s956 : std_logic_vector(33 downto 0) := (others => '0');
signal s957 : std_logic_vector(33 downto 0) := (others => '0');
signal s958 : std_logic_vector(33 downto 0) := (others => '0');
signal s959 : std_logic_vector(33 downto 0) := (others => '0');
signal s960 : std_logic_vector(33 downto 0) := (others => '0');
signal s961 : std_logic_vector(33 downto 0) := (others => '0');
signal s962 : std_logic_vector(33 downto 0) := (others => '0');
signal s963 : std_logic_vector(33 downto 0) := (others => '0');
signal s964 : std_logic_vector(33 downto 0) := (others => '0');
signal s965 : std_logic_vector(33 downto 0) := (others => '0');
signal s966 : std_logic_vector(33 downto 0) := (others => '0');
signal s967 : std_logic_vector(33 downto 0) := (others => '0');
signal s968 : std_logic_vector(33 downto 0) := (others => '0');
signal s969 : std_logic_vector(33 downto 0) := (others => '0');
signal s970 : std_logic_vector(33 downto 0) := (others => '0');
signal s971 : std_logic_vector(33 downto 0) := (others => '0');
signal s972 : std_logic_vector(33 downto 0) := (others => '0');
signal s973 : std_logic_vector(33 downto 0) := (others => '0');
signal s974 : std_logic_vector(33 downto 0) := (others => '0');
signal s975 : std_logic_vector(33 downto 0) := (others => '0');
signal s976 : std_logic_vector(33 downto 0) := (others => '0');
signal s977 : std_logic_vector(33 downto 0) := (others => '0');
signal s978 : std_logic_vector(33 downto 0) := (others => '0');
signal s979 : std_logic_vector(33 downto 0) := (others => '0');
signal s980 : std_logic_vector(33 downto 0) := (others => '0');
signal s981 : std_logic_vector(33 downto 0) := (others => '0');
signal s982 : std_logic_vector(33 downto 0) := (others => '0');
signal s983 : std_logic_vector(33 downto 0) := (others => '0');
signal s984 : std_logic_vector(33 downto 0) := (others => '0');
signal s985 : std_logic_vector(33 downto 0) := (others => '0');
signal s986 : std_logic_vector(33 downto 0) := (others => '0');
signal s987 : std_logic_vector(33 downto 0) := (others => '0');
signal s988 : std_logic_vector(33 downto 0) := (others => '0');
signal s989 : std_logic_vector(33 downto 0) := (others => '0');
signal s990 : std_logic_vector(33 downto 0) := (others => '0');
signal s991 : std_logic_vector(33 downto 0) := (others => '0');
signal s992 : std_logic_vector(33 downto 0) := (others => '0');
signal s993 : std_logic_vector(33 downto 0) := (others => '0');
signal s994 : std_logic_vector(33 downto 0) := (others => '0');
signal s995 : std_logic_vector(33 downto 0) := (others => '0');
signal s996 : std_logic_vector(33 downto 0) := (others => '0');
signal s997 : std_logic_vector(33 downto 0) := (others => '0');
signal s998 : std_logic_vector(33 downto 0) := (others => '0');
signal s999 : std_logic_vector(33 downto 0) := (others => '0');
signal s1000 : std_logic_vector(33 downto 0) := (others => '0');
signal s1001 : std_logic_vector(33 downto 0) := (others => '0');
signal s1002 : std_logic_vector(33 downto 0) := (others => '0');
signal s1003 : std_logic_vector(33 downto 0) := (others => '0');
signal s1004 : std_logic_vector(33 downto 0) := (others => '0');
signal s1005 : std_logic_vector(33 downto 0) := (others => '0');
signal s1006 : std_logic_vector(33 downto 0) := (others => '0');
signal s1007 : std_logic_vector(33 downto 0) := (others => '0');
signal s1008 : std_logic_vector(33 downto 0) := (others => '0');
signal s1009 : std_logic_vector(33 downto 0) := (others => '0');
signal s1010 : std_logic_vector(33 downto 0) := (others => '0');
signal s1011 : std_logic_vector(33 downto 0) := (others => '0');
signal s1012 : std_logic_vector(33 downto 0) := (others => '0');
signal s1013 : std_logic_vector(33 downto 0) := (others => '0');
signal s1014 : std_logic_vector(33 downto 0) := (others => '0');
signal s1015 : std_logic_vector(33 downto 0) := (others => '0');
signal s1016 : std_logic_vector(33 downto 0) := (others => '0');
signal s1017 : std_logic_vector(33 downto 0) := (others => '0');
signal s1018 : std_logic_vector(33 downto 0) := (others => '0');
signal s1019 : std_logic_vector(33 downto 0) := (others => '0');
signal s1020 : std_logic_vector(33 downto 0) := (others => '0');
signal s1021 : std_logic_vector(33 downto 0) := (others => '0');
signal s1022 : std_logic_vector(33 downto 0) := (others => '0');
signal s1023 : std_logic_vector(33 downto 0) := (others => '0');
signal s1024 : std_logic_vector(33 downto 0) := (others => '0');
signal s1025 : std_logic_vector(33 downto 0) := (others => '0');
signal s1026 : std_logic_vector(33 downto 0) := (others => '0');
signal s1027 : std_logic_vector(33 downto 0) := (others => '0');
signal s1028 : std_logic_vector(33 downto 0) := (others => '0');
signal s1029 : std_logic_vector(33 downto 0) := (others => '0');
signal s1030 : std_logic_vector(33 downto 0) := (others => '0');
signal s1031 : std_logic_vector(33 downto 0) := (others => '0');
signal s1032 : std_logic_vector(33 downto 0) := (others => '0');
signal s1033 : std_logic_vector(33 downto 0) := (others => '0');
signal s1034 : std_logic_vector(33 downto 0) := (others => '0');
signal s1035 : std_logic_vector(33 downto 0) := (others => '0');
signal s1036 : std_logic_vector(33 downto 0) := (others => '0');
signal s1037 : std_logic_vector(33 downto 0) := (others => '0');
signal s1038 : std_logic_vector(33 downto 0) := (others => '0');
signal s1039 : std_logic_vector(33 downto 0) := (others => '0');
signal s1040 : std_logic_vector(33 downto 0) := (others => '0');
signal s1041 : std_logic_vector(33 downto 0) := (others => '0');
signal s1042 : std_logic_vector(33 downto 0) := (others => '0');
signal s1043 : std_logic_vector(33 downto 0) := (others => '0');
signal s1044 : std_logic_vector(33 downto 0) := (others => '0');
signal s1045 : std_logic_vector(33 downto 0) := (others => '0');
signal s1046 : std_logic_vector(33 downto 0) := (others => '0');
signal s1047 : std_logic_vector(33 downto 0) := (others => '0');
signal s1048 : std_logic_vector(33 downto 0) := (others => '0');
signal s1049 : std_logic_vector(33 downto 0) := (others => '0');
signal s1050 : std_logic_vector(33 downto 0) := (others => '0');
signal s1051 : std_logic_vector(33 downto 0) := (others => '0');
signal s1052 : std_logic_vector(33 downto 0) := (others => '0');
signal s1053 : std_logic_vector(33 downto 0) := (others => '0');
signal s1054 : std_logic_vector(33 downto 0) := (others => '0');
signal s1055 : std_logic_vector(33 downto 0) := (others => '0');
signal s1056 : std_logic_vector(33 downto 0) := (others => '0');
signal s1057 : std_logic_vector(33 downto 0) := (others => '0');
signal s1058 : std_logic_vector(33 downto 0) := (others => '0');
signal s1059 : std_logic_vector(33 downto 0) := (others => '0');
signal s1060 : std_logic_vector(33 downto 0) := (others => '0');
signal s1061 : std_logic_vector(33 downto 0) := (others => '0');
signal s1062 : std_logic_vector(33 downto 0) := (others => '0');
signal s1063 : std_logic_vector(33 downto 0) := (others => '0');
signal s1064 : std_logic_vector(33 downto 0) := (others => '0');
signal s1065 : std_logic_vector(33 downto 0) := (others => '0');
signal s1066 : std_logic_vector(33 downto 0) := (others => '0');
signal s1067 : std_logic_vector(33 downto 0) := (others => '0');
signal s1068 : std_logic_vector(33 downto 0) := (others => '0');
signal s1069 : std_logic_vector(33 downto 0) := (others => '0');
signal s1070 : std_logic_vector(33 downto 0) := (others => '0');
signal s1071 : std_logic_vector(33 downto 0) := (others => '0');
signal s1072 : std_logic_vector(33 downto 0) := (others => '0');
signal s1073 : std_logic_vector(33 downto 0) := (others => '0');
signal s1074 : std_logic_vector(33 downto 0) := (others => '0');
signal s1075 : std_logic_vector(33 downto 0) := (others => '0');
signal s1076 : std_logic_vector(33 downto 0) := (others => '0');
signal s1077 : std_logic_vector(33 downto 0) := (others => '0');
signal s1078 : std_logic_vector(33 downto 0) := (others => '0');
signal s1079 : std_logic_vector(33 downto 0) := (others => '0');
signal s1080 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
      s558 <= "0000000000000000000000000000000000";
      s559 <= "0000000000000000000000000000000000";
      s560 <= "0000000000000000000000000000000000";
      s561 <= "0000000000000000000000000000000000";
      s562 <= "0000000000000000000000000000000000";
      s563 <= "0000000000000000000000000000000000";
      s564 <= "0000000000000000000000000000000000";
      s565 <= "0000000000000000000000000000000000";
      s566 <= "0000000000000000000000000000000000";
      s567 <= "0000000000000000000000000000000000";
      s568 <= "0000000000000000000000000000000000";
      s569 <= "0000000000000000000000000000000000";
      s570 <= "0000000000000000000000000000000000";
      s571 <= "0000000000000000000000000000000000";
      s572 <= "0000000000000000000000000000000000";
      s573 <= "0000000000000000000000000000000000";
      s574 <= "0000000000000000000000000000000000";
      s575 <= "0000000000000000000000000000000000";
      s576 <= "0000000000000000000000000000000000";
      s577 <= "0000000000000000000000000000000000";
      s578 <= "0000000000000000000000000000000000";
      s579 <= "0000000000000000000000000000000000";
      s580 <= "0000000000000000000000000000000000";
      s581 <= "0000000000000000000000000000000000";
      s582 <= "0000000000000000000000000000000000";
      s583 <= "0000000000000000000000000000000000";
      s584 <= "0000000000000000000000000000000000";
      s585 <= "0000000000000000000000000000000000";
      s586 <= "0000000000000000000000000000000000";
      s587 <= "0000000000000000000000000000000000";
      s588 <= "0000000000000000000000000000000000";
      s589 <= "0000000000000000000000000000000000";
      s590 <= "0000000000000000000000000000000000";
      s591 <= "0000000000000000000000000000000000";
      s592 <= "0000000000000000000000000000000000";
      s593 <= "0000000000000000000000000000000000";
      s594 <= "0000000000000000000000000000000000";
      s595 <= "0000000000000000000000000000000000";
      s596 <= "0000000000000000000000000000000000";
      s597 <= "0000000000000000000000000000000000";
      s598 <= "0000000000000000000000000000000000";
      s599 <= "0000000000000000000000000000000000";
      s600 <= "0000000000000000000000000000000000";
      s601 <= "0000000000000000000000000000000000";
      s602 <= "0000000000000000000000000000000000";
      s603 <= "0000000000000000000000000000000000";
      s604 <= "0000000000000000000000000000000000";
      s605 <= "0000000000000000000000000000000000";
      s606 <= "0000000000000000000000000000000000";
      s607 <= "0000000000000000000000000000000000";
      s608 <= "0000000000000000000000000000000000";
      s609 <= "0000000000000000000000000000000000";
      s610 <= "0000000000000000000000000000000000";
      s611 <= "0000000000000000000000000000000000";
      s612 <= "0000000000000000000000000000000000";
      s613 <= "0000000000000000000000000000000000";
      s614 <= "0000000000000000000000000000000000";
      s615 <= "0000000000000000000000000000000000";
      s616 <= "0000000000000000000000000000000000";
      s617 <= "0000000000000000000000000000000000";
      s618 <= "0000000000000000000000000000000000";
      s619 <= "0000000000000000000000000000000000";
      s620 <= "0000000000000000000000000000000000";
      s621 <= "0000000000000000000000000000000000";
      s622 <= "0000000000000000000000000000000000";
      s623 <= "0000000000000000000000000000000000";
      s624 <= "0000000000000000000000000000000000";
      s625 <= "0000000000000000000000000000000000";
      s626 <= "0000000000000000000000000000000000";
      s627 <= "0000000000000000000000000000000000";
      s628 <= "0000000000000000000000000000000000";
      s629 <= "0000000000000000000000000000000000";
      s630 <= "0000000000000000000000000000000000";
      s631 <= "0000000000000000000000000000000000";
      s632 <= "0000000000000000000000000000000000";
      s633 <= "0000000000000000000000000000000000";
      s634 <= "0000000000000000000000000000000000";
      s635 <= "0000000000000000000000000000000000";
      s636 <= "0000000000000000000000000000000000";
      s637 <= "0000000000000000000000000000000000";
      s638 <= "0000000000000000000000000000000000";
      s639 <= "0000000000000000000000000000000000";
      s640 <= "0000000000000000000000000000000000";
      s641 <= "0000000000000000000000000000000000";
      s642 <= "0000000000000000000000000000000000";
      s643 <= "0000000000000000000000000000000000";
      s644 <= "0000000000000000000000000000000000";
      s645 <= "0000000000000000000000000000000000";
      s646 <= "0000000000000000000000000000000000";
      s647 <= "0000000000000000000000000000000000";
      s648 <= "0000000000000000000000000000000000";
      s649 <= "0000000000000000000000000000000000";
      s650 <= "0000000000000000000000000000000000";
      s651 <= "0000000000000000000000000000000000";
      s652 <= "0000000000000000000000000000000000";
      s653 <= "0000000000000000000000000000000000";
      s654 <= "0000000000000000000000000000000000";
      s655 <= "0000000000000000000000000000000000";
      s656 <= "0000000000000000000000000000000000";
      s657 <= "0000000000000000000000000000000000";
      s658 <= "0000000000000000000000000000000000";
      s659 <= "0000000000000000000000000000000000";
      s660 <= "0000000000000000000000000000000000";
      s661 <= "0000000000000000000000000000000000";
      s662 <= "0000000000000000000000000000000000";
      s663 <= "0000000000000000000000000000000000";
      s664 <= "0000000000000000000000000000000000";
      s665 <= "0000000000000000000000000000000000";
      s666 <= "0000000000000000000000000000000000";
      s667 <= "0000000000000000000000000000000000";
      s668 <= "0000000000000000000000000000000000";
      s669 <= "0000000000000000000000000000000000";
      s670 <= "0000000000000000000000000000000000";
      s671 <= "0000000000000000000000000000000000";
      s672 <= "0000000000000000000000000000000000";
      s673 <= "0000000000000000000000000000000000";
      s674 <= "0000000000000000000000000000000000";
      s675 <= "0000000000000000000000000000000000";
      s676 <= "0000000000000000000000000000000000";
      s677 <= "0000000000000000000000000000000000";
      s678 <= "0000000000000000000000000000000000";
      s679 <= "0000000000000000000000000000000000";
      s680 <= "0000000000000000000000000000000000";
      s681 <= "0000000000000000000000000000000000";
      s682 <= "0000000000000000000000000000000000";
      s683 <= "0000000000000000000000000000000000";
      s684 <= "0000000000000000000000000000000000";
      s685 <= "0000000000000000000000000000000000";
      s686 <= "0000000000000000000000000000000000";
      s687 <= "0000000000000000000000000000000000";
      s688 <= "0000000000000000000000000000000000";
      s689 <= "0000000000000000000000000000000000";
      s690 <= "0000000000000000000000000000000000";
      s691 <= "0000000000000000000000000000000000";
      s692 <= "0000000000000000000000000000000000";
      s693 <= "0000000000000000000000000000000000";
      s694 <= "0000000000000000000000000000000000";
      s695 <= "0000000000000000000000000000000000";
      s696 <= "0000000000000000000000000000000000";
      s697 <= "0000000000000000000000000000000000";
      s698 <= "0000000000000000000000000000000000";
      s699 <= "0000000000000000000000000000000000";
      s700 <= "0000000000000000000000000000000000";
      s701 <= "0000000000000000000000000000000000";
      s702 <= "0000000000000000000000000000000000";
      s703 <= "0000000000000000000000000000000000";
      s704 <= "0000000000000000000000000000000000";
      s705 <= "0000000000000000000000000000000000";
      s706 <= "0000000000000000000000000000000000";
      s707 <= "0000000000000000000000000000000000";
      s708 <= "0000000000000000000000000000000000";
      s709 <= "0000000000000000000000000000000000";
      s710 <= "0000000000000000000000000000000000";
      s711 <= "0000000000000000000000000000000000";
      s712 <= "0000000000000000000000000000000000";
      s713 <= "0000000000000000000000000000000000";
      s714 <= "0000000000000000000000000000000000";
      s715 <= "0000000000000000000000000000000000";
      s716 <= "0000000000000000000000000000000000";
      s717 <= "0000000000000000000000000000000000";
      s718 <= "0000000000000000000000000000000000";
      s719 <= "0000000000000000000000000000000000";
      s720 <= "0000000000000000000000000000000000";
      s721 <= "0000000000000000000000000000000000";
      s722 <= "0000000000000000000000000000000000";
      s723 <= "0000000000000000000000000000000000";
      s724 <= "0000000000000000000000000000000000";
      s725 <= "0000000000000000000000000000000000";
      s726 <= "0000000000000000000000000000000000";
      s727 <= "0000000000000000000000000000000000";
      s728 <= "0000000000000000000000000000000000";
      s729 <= "0000000000000000000000000000000000";
      s730 <= "0000000000000000000000000000000000";
      s731 <= "0000000000000000000000000000000000";
      s732 <= "0000000000000000000000000000000000";
      s733 <= "0000000000000000000000000000000000";
      s734 <= "0000000000000000000000000000000000";
      s735 <= "0000000000000000000000000000000000";
      s736 <= "0000000000000000000000000000000000";
      s737 <= "0000000000000000000000000000000000";
      s738 <= "0000000000000000000000000000000000";
      s739 <= "0000000000000000000000000000000000";
      s740 <= "0000000000000000000000000000000000";
      s741 <= "0000000000000000000000000000000000";
      s742 <= "0000000000000000000000000000000000";
      s743 <= "0000000000000000000000000000000000";
      s744 <= "0000000000000000000000000000000000";
      s745 <= "0000000000000000000000000000000000";
      s746 <= "0000000000000000000000000000000000";
      s747 <= "0000000000000000000000000000000000";
      s748 <= "0000000000000000000000000000000000";
      s749 <= "0000000000000000000000000000000000";
      s750 <= "0000000000000000000000000000000000";
      s751 <= "0000000000000000000000000000000000";
      s752 <= "0000000000000000000000000000000000";
      s753 <= "0000000000000000000000000000000000";
      s754 <= "0000000000000000000000000000000000";
      s755 <= "0000000000000000000000000000000000";
      s756 <= "0000000000000000000000000000000000";
      s757 <= "0000000000000000000000000000000000";
      s758 <= "0000000000000000000000000000000000";
      s759 <= "0000000000000000000000000000000000";
      s760 <= "0000000000000000000000000000000000";
      s761 <= "0000000000000000000000000000000000";
      s762 <= "0000000000000000000000000000000000";
      s763 <= "0000000000000000000000000000000000";
      s764 <= "0000000000000000000000000000000000";
      s765 <= "0000000000000000000000000000000000";
      s766 <= "0000000000000000000000000000000000";
      s767 <= "0000000000000000000000000000000000";
      s768 <= "0000000000000000000000000000000000";
      s769 <= "0000000000000000000000000000000000";
      s770 <= "0000000000000000000000000000000000";
      s771 <= "0000000000000000000000000000000000";
      s772 <= "0000000000000000000000000000000000";
      s773 <= "0000000000000000000000000000000000";
      s774 <= "0000000000000000000000000000000000";
      s775 <= "0000000000000000000000000000000000";
      s776 <= "0000000000000000000000000000000000";
      s777 <= "0000000000000000000000000000000000";
      s778 <= "0000000000000000000000000000000000";
      s779 <= "0000000000000000000000000000000000";
      s780 <= "0000000000000000000000000000000000";
      s781 <= "0000000000000000000000000000000000";
      s782 <= "0000000000000000000000000000000000";
      s783 <= "0000000000000000000000000000000000";
      s784 <= "0000000000000000000000000000000000";
      s785 <= "0000000000000000000000000000000000";
      s786 <= "0000000000000000000000000000000000";
      s787 <= "0000000000000000000000000000000000";
      s788 <= "0000000000000000000000000000000000";
      s789 <= "0000000000000000000000000000000000";
      s790 <= "0000000000000000000000000000000000";
      s791 <= "0000000000000000000000000000000000";
      s792 <= "0000000000000000000000000000000000";
      s793 <= "0000000000000000000000000000000000";
      s794 <= "0000000000000000000000000000000000";
      s795 <= "0000000000000000000000000000000000";
      s796 <= "0000000000000000000000000000000000";
      s797 <= "0000000000000000000000000000000000";
      s798 <= "0000000000000000000000000000000000";
      s799 <= "0000000000000000000000000000000000";
      s800 <= "0000000000000000000000000000000000";
      s801 <= "0000000000000000000000000000000000";
      s802 <= "0000000000000000000000000000000000";
      s803 <= "0000000000000000000000000000000000";
      s804 <= "0000000000000000000000000000000000";
      s805 <= "0000000000000000000000000000000000";
      s806 <= "0000000000000000000000000000000000";
      s807 <= "0000000000000000000000000000000000";
      s808 <= "0000000000000000000000000000000000";
      s809 <= "0000000000000000000000000000000000";
      s810 <= "0000000000000000000000000000000000";
      s811 <= "0000000000000000000000000000000000";
      s812 <= "0000000000000000000000000000000000";
      s813 <= "0000000000000000000000000000000000";
      s814 <= "0000000000000000000000000000000000";
      s815 <= "0000000000000000000000000000000000";
      s816 <= "0000000000000000000000000000000000";
      s817 <= "0000000000000000000000000000000000";
      s818 <= "0000000000000000000000000000000000";
      s819 <= "0000000000000000000000000000000000";
      s820 <= "0000000000000000000000000000000000";
      s821 <= "0000000000000000000000000000000000";
      s822 <= "0000000000000000000000000000000000";
      s823 <= "0000000000000000000000000000000000";
      s824 <= "0000000000000000000000000000000000";
      s825 <= "0000000000000000000000000000000000";
      s826 <= "0000000000000000000000000000000000";
      s827 <= "0000000000000000000000000000000000";
      s828 <= "0000000000000000000000000000000000";
      s829 <= "0000000000000000000000000000000000";
      s830 <= "0000000000000000000000000000000000";
      s831 <= "0000000000000000000000000000000000";
      s832 <= "0000000000000000000000000000000000";
      s833 <= "0000000000000000000000000000000000";
      s834 <= "0000000000000000000000000000000000";
      s835 <= "0000000000000000000000000000000000";
      s836 <= "0000000000000000000000000000000000";
      s837 <= "0000000000000000000000000000000000";
      s838 <= "0000000000000000000000000000000000";
      s839 <= "0000000000000000000000000000000000";
      s840 <= "0000000000000000000000000000000000";
      s841 <= "0000000000000000000000000000000000";
      s842 <= "0000000000000000000000000000000000";
      s843 <= "0000000000000000000000000000000000";
      s844 <= "0000000000000000000000000000000000";
      s845 <= "0000000000000000000000000000000000";
      s846 <= "0000000000000000000000000000000000";
      s847 <= "0000000000000000000000000000000000";
      s848 <= "0000000000000000000000000000000000";
      s849 <= "0000000000000000000000000000000000";
      s850 <= "0000000000000000000000000000000000";
      s851 <= "0000000000000000000000000000000000";
      s852 <= "0000000000000000000000000000000000";
      s853 <= "0000000000000000000000000000000000";
      s854 <= "0000000000000000000000000000000000";
      s855 <= "0000000000000000000000000000000000";
      s856 <= "0000000000000000000000000000000000";
      s857 <= "0000000000000000000000000000000000";
      s858 <= "0000000000000000000000000000000000";
      s859 <= "0000000000000000000000000000000000";
      s860 <= "0000000000000000000000000000000000";
      s861 <= "0000000000000000000000000000000000";
      s862 <= "0000000000000000000000000000000000";
      s863 <= "0000000000000000000000000000000000";
      s864 <= "0000000000000000000000000000000000";
      s865 <= "0000000000000000000000000000000000";
      s866 <= "0000000000000000000000000000000000";
      s867 <= "0000000000000000000000000000000000";
      s868 <= "0000000000000000000000000000000000";
      s869 <= "0000000000000000000000000000000000";
      s870 <= "0000000000000000000000000000000000";
      s871 <= "0000000000000000000000000000000000";
      s872 <= "0000000000000000000000000000000000";
      s873 <= "0000000000000000000000000000000000";
      s874 <= "0000000000000000000000000000000000";
      s875 <= "0000000000000000000000000000000000";
      s876 <= "0000000000000000000000000000000000";
      s877 <= "0000000000000000000000000000000000";
      s878 <= "0000000000000000000000000000000000";
      s879 <= "0000000000000000000000000000000000";
      s880 <= "0000000000000000000000000000000000";
      s881 <= "0000000000000000000000000000000000";
      s882 <= "0000000000000000000000000000000000";
      s883 <= "0000000000000000000000000000000000";
      s884 <= "0000000000000000000000000000000000";
      s885 <= "0000000000000000000000000000000000";
      s886 <= "0000000000000000000000000000000000";
      s887 <= "0000000000000000000000000000000000";
      s888 <= "0000000000000000000000000000000000";
      s889 <= "0000000000000000000000000000000000";
      s890 <= "0000000000000000000000000000000000";
      s891 <= "0000000000000000000000000000000000";
      s892 <= "0000000000000000000000000000000000";
      s893 <= "0000000000000000000000000000000000";
      s894 <= "0000000000000000000000000000000000";
      s895 <= "0000000000000000000000000000000000";
      s896 <= "0000000000000000000000000000000000";
      s897 <= "0000000000000000000000000000000000";
      s898 <= "0000000000000000000000000000000000";
      s899 <= "0000000000000000000000000000000000";
      s900 <= "0000000000000000000000000000000000";
      s901 <= "0000000000000000000000000000000000";
      s902 <= "0000000000000000000000000000000000";
      s903 <= "0000000000000000000000000000000000";
      s904 <= "0000000000000000000000000000000000";
      s905 <= "0000000000000000000000000000000000";
      s906 <= "0000000000000000000000000000000000";
      s907 <= "0000000000000000000000000000000000";
      s908 <= "0000000000000000000000000000000000";
      s909 <= "0000000000000000000000000000000000";
      s910 <= "0000000000000000000000000000000000";
      s911 <= "0000000000000000000000000000000000";
      s912 <= "0000000000000000000000000000000000";
      s913 <= "0000000000000000000000000000000000";
      s914 <= "0000000000000000000000000000000000";
      s915 <= "0000000000000000000000000000000000";
      s916 <= "0000000000000000000000000000000000";
      s917 <= "0000000000000000000000000000000000";
      s918 <= "0000000000000000000000000000000000";
      s919 <= "0000000000000000000000000000000000";
      s920 <= "0000000000000000000000000000000000";
      s921 <= "0000000000000000000000000000000000";
      s922 <= "0000000000000000000000000000000000";
      s923 <= "0000000000000000000000000000000000";
      s924 <= "0000000000000000000000000000000000";
      s925 <= "0000000000000000000000000000000000";
      s926 <= "0000000000000000000000000000000000";
      s927 <= "0000000000000000000000000000000000";
      s928 <= "0000000000000000000000000000000000";
      s929 <= "0000000000000000000000000000000000";
      s930 <= "0000000000000000000000000000000000";
      s931 <= "0000000000000000000000000000000000";
      s932 <= "0000000000000000000000000000000000";
      s933 <= "0000000000000000000000000000000000";
      s934 <= "0000000000000000000000000000000000";
      s935 <= "0000000000000000000000000000000000";
      s936 <= "0000000000000000000000000000000000";
      s937 <= "0000000000000000000000000000000000";
      s938 <= "0000000000000000000000000000000000";
      s939 <= "0000000000000000000000000000000000";
      s940 <= "0000000000000000000000000000000000";
      s941 <= "0000000000000000000000000000000000";
      s942 <= "0000000000000000000000000000000000";
      s943 <= "0000000000000000000000000000000000";
      s944 <= "0000000000000000000000000000000000";
      s945 <= "0000000000000000000000000000000000";
      s946 <= "0000000000000000000000000000000000";
      s947 <= "0000000000000000000000000000000000";
      s948 <= "0000000000000000000000000000000000";
      s949 <= "0000000000000000000000000000000000";
      s950 <= "0000000000000000000000000000000000";
      s951 <= "0000000000000000000000000000000000";
      s952 <= "0000000000000000000000000000000000";
      s953 <= "0000000000000000000000000000000000";
      s954 <= "0000000000000000000000000000000000";
      s955 <= "0000000000000000000000000000000000";
      s956 <= "0000000000000000000000000000000000";
      s957 <= "0000000000000000000000000000000000";
      s958 <= "0000000000000000000000000000000000";
      s959 <= "0000000000000000000000000000000000";
      s960 <= "0000000000000000000000000000000000";
      s961 <= "0000000000000000000000000000000000";
      s962 <= "0000000000000000000000000000000000";
      s963 <= "0000000000000000000000000000000000";
      s964 <= "0000000000000000000000000000000000";
      s965 <= "0000000000000000000000000000000000";
      s966 <= "0000000000000000000000000000000000";
      s967 <= "0000000000000000000000000000000000";
      s968 <= "0000000000000000000000000000000000";
      s969 <= "0000000000000000000000000000000000";
      s970 <= "0000000000000000000000000000000000";
      s971 <= "0000000000000000000000000000000000";
      s972 <= "0000000000000000000000000000000000";
      s973 <= "0000000000000000000000000000000000";
      s974 <= "0000000000000000000000000000000000";
      s975 <= "0000000000000000000000000000000000";
      s976 <= "0000000000000000000000000000000000";
      s977 <= "0000000000000000000000000000000000";
      s978 <= "0000000000000000000000000000000000";
      s979 <= "0000000000000000000000000000000000";
      s980 <= "0000000000000000000000000000000000";
      s981 <= "0000000000000000000000000000000000";
      s982 <= "0000000000000000000000000000000000";
      s983 <= "0000000000000000000000000000000000";
      s984 <= "0000000000000000000000000000000000";
      s985 <= "0000000000000000000000000000000000";
      s986 <= "0000000000000000000000000000000000";
      s987 <= "0000000000000000000000000000000000";
      s988 <= "0000000000000000000000000000000000";
      s989 <= "0000000000000000000000000000000000";
      s990 <= "0000000000000000000000000000000000";
      s991 <= "0000000000000000000000000000000000";
      s992 <= "0000000000000000000000000000000000";
      s993 <= "0000000000000000000000000000000000";
      s994 <= "0000000000000000000000000000000000";
      s995 <= "0000000000000000000000000000000000";
      s996 <= "0000000000000000000000000000000000";
      s997 <= "0000000000000000000000000000000000";
      s998 <= "0000000000000000000000000000000000";
      s999 <= "0000000000000000000000000000000000";
      s1000 <= "0000000000000000000000000000000000";
      s1001 <= "0000000000000000000000000000000000";
      s1002 <= "0000000000000000000000000000000000";
      s1003 <= "0000000000000000000000000000000000";
      s1004 <= "0000000000000000000000000000000000";
      s1005 <= "0000000000000000000000000000000000";
      s1006 <= "0000000000000000000000000000000000";
      s1007 <= "0000000000000000000000000000000000";
      s1008 <= "0000000000000000000000000000000000";
      s1009 <= "0000000000000000000000000000000000";
      s1010 <= "0000000000000000000000000000000000";
      s1011 <= "0000000000000000000000000000000000";
      s1012 <= "0000000000000000000000000000000000";
      s1013 <= "0000000000000000000000000000000000";
      s1014 <= "0000000000000000000000000000000000";
      s1015 <= "0000000000000000000000000000000000";
      s1016 <= "0000000000000000000000000000000000";
      s1017 <= "0000000000000000000000000000000000";
      s1018 <= "0000000000000000000000000000000000";
      s1019 <= "0000000000000000000000000000000000";
      s1020 <= "0000000000000000000000000000000000";
      s1021 <= "0000000000000000000000000000000000";
      s1022 <= "0000000000000000000000000000000000";
      s1023 <= "0000000000000000000000000000000000";
      s1024 <= "0000000000000000000000000000000000";
      s1025 <= "0000000000000000000000000000000000";
      s1026 <= "0000000000000000000000000000000000";
      s1027 <= "0000000000000000000000000000000000";
      s1028 <= "0000000000000000000000000000000000";
      s1029 <= "0000000000000000000000000000000000";
      s1030 <= "0000000000000000000000000000000000";
      s1031 <= "0000000000000000000000000000000000";
      s1032 <= "0000000000000000000000000000000000";
      s1033 <= "0000000000000000000000000000000000";
      s1034 <= "0000000000000000000000000000000000";
      s1035 <= "0000000000000000000000000000000000";
      s1036 <= "0000000000000000000000000000000000";
      s1037 <= "0000000000000000000000000000000000";
      s1038 <= "0000000000000000000000000000000000";
      s1039 <= "0000000000000000000000000000000000";
      s1040 <= "0000000000000000000000000000000000";
      s1041 <= "0000000000000000000000000000000000";
      s1042 <= "0000000000000000000000000000000000";
      s1043 <= "0000000000000000000000000000000000";
      s1044 <= "0000000000000000000000000000000000";
      s1045 <= "0000000000000000000000000000000000";
      s1046 <= "0000000000000000000000000000000000";
      s1047 <= "0000000000000000000000000000000000";
      s1048 <= "0000000000000000000000000000000000";
      s1049 <= "0000000000000000000000000000000000";
      s1050 <= "0000000000000000000000000000000000";
      s1051 <= "0000000000000000000000000000000000";
      s1052 <= "0000000000000000000000000000000000";
      s1053 <= "0000000000000000000000000000000000";
      s1054 <= "0000000000000000000000000000000000";
      s1055 <= "0000000000000000000000000000000000";
      s1056 <= "0000000000000000000000000000000000";
      s1057 <= "0000000000000000000000000000000000";
      s1058 <= "0000000000000000000000000000000000";
      s1059 <= "0000000000000000000000000000000000";
      s1060 <= "0000000000000000000000000000000000";
      s1061 <= "0000000000000000000000000000000000";
      s1062 <= "0000000000000000000000000000000000";
      s1063 <= "0000000000000000000000000000000000";
      s1064 <= "0000000000000000000000000000000000";
      s1065 <= "0000000000000000000000000000000000";
      s1066 <= "0000000000000000000000000000000000";
      s1067 <= "0000000000000000000000000000000000";
      s1068 <= "0000000000000000000000000000000000";
      s1069 <= "0000000000000000000000000000000000";
      s1070 <= "0000000000000000000000000000000000";
      s1071 <= "0000000000000000000000000000000000";
      s1072 <= "0000000000000000000000000000000000";
      s1073 <= "0000000000000000000000000000000000";
      s1074 <= "0000000000000000000000000000000000";
      s1075 <= "0000000000000000000000000000000000";
      s1076 <= "0000000000000000000000000000000000";
      s1077 <= "0000000000000000000000000000000000";
      s1078 <= "0000000000000000000000000000000000";
      s1079 <= "0000000000000000000000000000000000";
      s1080 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      s558 <= s557;
      s559 <= s558;
      s560 <= s559;
      s561 <= s560;
      s562 <= s561;
      s563 <= s562;
      s564 <= s563;
      s565 <= s564;
      s566 <= s565;
      s567 <= s566;
      s568 <= s567;
      s569 <= s568;
      s570 <= s569;
      s571 <= s570;
      s572 <= s571;
      s573 <= s572;
      s574 <= s573;
      s575 <= s574;
      s576 <= s575;
      s577 <= s576;
      s578 <= s577;
      s579 <= s578;
      s580 <= s579;
      s581 <= s580;
      s582 <= s581;
      s583 <= s582;
      s584 <= s583;
      s585 <= s584;
      s586 <= s585;
      s587 <= s586;
      s588 <= s587;
      s589 <= s588;
      s590 <= s589;
      s591 <= s590;
      s592 <= s591;
      s593 <= s592;
      s594 <= s593;
      s595 <= s594;
      s596 <= s595;
      s597 <= s596;
      s598 <= s597;
      s599 <= s598;
      s600 <= s599;
      s601 <= s600;
      s602 <= s601;
      s603 <= s602;
      s604 <= s603;
      s605 <= s604;
      s606 <= s605;
      s607 <= s606;
      s608 <= s607;
      s609 <= s608;
      s610 <= s609;
      s611 <= s610;
      s612 <= s611;
      s613 <= s612;
      s614 <= s613;
      s615 <= s614;
      s616 <= s615;
      s617 <= s616;
      s618 <= s617;
      s619 <= s618;
      s620 <= s619;
      s621 <= s620;
      s622 <= s621;
      s623 <= s622;
      s624 <= s623;
      s625 <= s624;
      s626 <= s625;
      s627 <= s626;
      s628 <= s627;
      s629 <= s628;
      s630 <= s629;
      s631 <= s630;
      s632 <= s631;
      s633 <= s632;
      s634 <= s633;
      s635 <= s634;
      s636 <= s635;
      s637 <= s636;
      s638 <= s637;
      s639 <= s638;
      s640 <= s639;
      s641 <= s640;
      s642 <= s641;
      s643 <= s642;
      s644 <= s643;
      s645 <= s644;
      s646 <= s645;
      s647 <= s646;
      s648 <= s647;
      s649 <= s648;
      s650 <= s649;
      s651 <= s650;
      s652 <= s651;
      s653 <= s652;
      s654 <= s653;
      s655 <= s654;
      s656 <= s655;
      s657 <= s656;
      s658 <= s657;
      s659 <= s658;
      s660 <= s659;
      s661 <= s660;
      s662 <= s661;
      s663 <= s662;
      s664 <= s663;
      s665 <= s664;
      s666 <= s665;
      s667 <= s666;
      s668 <= s667;
      s669 <= s668;
      s670 <= s669;
      s671 <= s670;
      s672 <= s671;
      s673 <= s672;
      s674 <= s673;
      s675 <= s674;
      s676 <= s675;
      s677 <= s676;
      s678 <= s677;
      s679 <= s678;
      s680 <= s679;
      s681 <= s680;
      s682 <= s681;
      s683 <= s682;
      s684 <= s683;
      s685 <= s684;
      s686 <= s685;
      s687 <= s686;
      s688 <= s687;
      s689 <= s688;
      s690 <= s689;
      s691 <= s690;
      s692 <= s691;
      s693 <= s692;
      s694 <= s693;
      s695 <= s694;
      s696 <= s695;
      s697 <= s696;
      s698 <= s697;
      s699 <= s698;
      s700 <= s699;
      s701 <= s700;
      s702 <= s701;
      s703 <= s702;
      s704 <= s703;
      s705 <= s704;
      s706 <= s705;
      s707 <= s706;
      s708 <= s707;
      s709 <= s708;
      s710 <= s709;
      s711 <= s710;
      s712 <= s711;
      s713 <= s712;
      s714 <= s713;
      s715 <= s714;
      s716 <= s715;
      s717 <= s716;
      s718 <= s717;
      s719 <= s718;
      s720 <= s719;
      s721 <= s720;
      s722 <= s721;
      s723 <= s722;
      s724 <= s723;
      s725 <= s724;
      s726 <= s725;
      s727 <= s726;
      s728 <= s727;
      s729 <= s728;
      s730 <= s729;
      s731 <= s730;
      s732 <= s731;
      s733 <= s732;
      s734 <= s733;
      s735 <= s734;
      s736 <= s735;
      s737 <= s736;
      s738 <= s737;
      s739 <= s738;
      s740 <= s739;
      s741 <= s740;
      s742 <= s741;
      s743 <= s742;
      s744 <= s743;
      s745 <= s744;
      s746 <= s745;
      s747 <= s746;
      s748 <= s747;
      s749 <= s748;
      s750 <= s749;
      s751 <= s750;
      s752 <= s751;
      s753 <= s752;
      s754 <= s753;
      s755 <= s754;
      s756 <= s755;
      s757 <= s756;
      s758 <= s757;
      s759 <= s758;
      s760 <= s759;
      s761 <= s760;
      s762 <= s761;
      s763 <= s762;
      s764 <= s763;
      s765 <= s764;
      s766 <= s765;
      s767 <= s766;
      s768 <= s767;
      s769 <= s768;
      s770 <= s769;
      s771 <= s770;
      s772 <= s771;
      s773 <= s772;
      s774 <= s773;
      s775 <= s774;
      s776 <= s775;
      s777 <= s776;
      s778 <= s777;
      s779 <= s778;
      s780 <= s779;
      s781 <= s780;
      s782 <= s781;
      s783 <= s782;
      s784 <= s783;
      s785 <= s784;
      s786 <= s785;
      s787 <= s786;
      s788 <= s787;
      s789 <= s788;
      s790 <= s789;
      s791 <= s790;
      s792 <= s791;
      s793 <= s792;
      s794 <= s793;
      s795 <= s794;
      s796 <= s795;
      s797 <= s796;
      s798 <= s797;
      s799 <= s798;
      s800 <= s799;
      s801 <= s800;
      s802 <= s801;
      s803 <= s802;
      s804 <= s803;
      s805 <= s804;
      s806 <= s805;
      s807 <= s806;
      s808 <= s807;
      s809 <= s808;
      s810 <= s809;
      s811 <= s810;
      s812 <= s811;
      s813 <= s812;
      s814 <= s813;
      s815 <= s814;
      s816 <= s815;
      s817 <= s816;
      s818 <= s817;
      s819 <= s818;
      s820 <= s819;
      s821 <= s820;
      s822 <= s821;
      s823 <= s822;
      s824 <= s823;
      s825 <= s824;
      s826 <= s825;
      s827 <= s826;
      s828 <= s827;
      s829 <= s828;
      s830 <= s829;
      s831 <= s830;
      s832 <= s831;
      s833 <= s832;
      s834 <= s833;
      s835 <= s834;
      s836 <= s835;
      s837 <= s836;
      s838 <= s837;
      s839 <= s838;
      s840 <= s839;
      s841 <= s840;
      s842 <= s841;
      s843 <= s842;
      s844 <= s843;
      s845 <= s844;
      s846 <= s845;
      s847 <= s846;
      s848 <= s847;
      s849 <= s848;
      s850 <= s849;
      s851 <= s850;
      s852 <= s851;
      s853 <= s852;
      s854 <= s853;
      s855 <= s854;
      s856 <= s855;
      s857 <= s856;
      s858 <= s857;
      s859 <= s858;
      s860 <= s859;
      s861 <= s860;
      s862 <= s861;
      s863 <= s862;
      s864 <= s863;
      s865 <= s864;
      s866 <= s865;
      s867 <= s866;
      s868 <= s867;
      s869 <= s868;
      s870 <= s869;
      s871 <= s870;
      s872 <= s871;
      s873 <= s872;
      s874 <= s873;
      s875 <= s874;
      s876 <= s875;
      s877 <= s876;
      s878 <= s877;
      s879 <= s878;
      s880 <= s879;
      s881 <= s880;
      s882 <= s881;
      s883 <= s882;
      s884 <= s883;
      s885 <= s884;
      s886 <= s885;
      s887 <= s886;
      s888 <= s887;
      s889 <= s888;
      s890 <= s889;
      s891 <= s890;
      s892 <= s891;
      s893 <= s892;
      s894 <= s893;
      s895 <= s894;
      s896 <= s895;
      s897 <= s896;
      s898 <= s897;
      s899 <= s898;
      s900 <= s899;
      s901 <= s900;
      s902 <= s901;
      s903 <= s902;
      s904 <= s903;
      s905 <= s904;
      s906 <= s905;
      s907 <= s906;
      s908 <= s907;
      s909 <= s908;
      s910 <= s909;
      s911 <= s910;
      s912 <= s911;
      s913 <= s912;
      s914 <= s913;
      s915 <= s914;
      s916 <= s915;
      s917 <= s916;
      s918 <= s917;
      s919 <= s918;
      s920 <= s919;
      s921 <= s920;
      s922 <= s921;
      s923 <= s922;
      s924 <= s923;
      s925 <= s924;
      s926 <= s925;
      s927 <= s926;
      s928 <= s927;
      s929 <= s928;
      s930 <= s929;
      s931 <= s930;
      s932 <= s931;
      s933 <= s932;
      s934 <= s933;
      s935 <= s934;
      s936 <= s935;
      s937 <= s936;
      s938 <= s937;
      s939 <= s938;
      s940 <= s939;
      s941 <= s940;
      s942 <= s941;
      s943 <= s942;
      s944 <= s943;
      s945 <= s944;
      s946 <= s945;
      s947 <= s946;
      s948 <= s947;
      s949 <= s948;
      s950 <= s949;
      s951 <= s950;
      s952 <= s951;
      s953 <= s952;
      s954 <= s953;
      s955 <= s954;
      s956 <= s955;
      s957 <= s956;
      s958 <= s957;
      s959 <= s958;
      s960 <= s959;
      s961 <= s960;
      s962 <= s961;
      s963 <= s962;
      s964 <= s963;
      s965 <= s964;
      s966 <= s965;
      s967 <= s966;
      s968 <= s967;
      s969 <= s968;
      s970 <= s969;
      s971 <= s970;
      s972 <= s971;
      s973 <= s972;
      s974 <= s973;
      s975 <= s974;
      s976 <= s975;
      s977 <= s976;
      s978 <= s977;
      s979 <= s978;
      s980 <= s979;
      s981 <= s980;
      s982 <= s981;
      s983 <= s982;
      s984 <= s983;
      s985 <= s984;
      s986 <= s985;
      s987 <= s986;
      s988 <= s987;
      s989 <= s988;
      s990 <= s989;
      s991 <= s990;
      s992 <= s991;
      s993 <= s992;
      s994 <= s993;
      s995 <= s994;
      s996 <= s995;
      s997 <= s996;
      s998 <= s997;
      s999 <= s998;
      s1000 <= s999;
      s1001 <= s1000;
      s1002 <= s1001;
      s1003 <= s1002;
      s1004 <= s1003;
      s1005 <= s1004;
      s1006 <= s1005;
      s1007 <= s1006;
      s1008 <= s1007;
      s1009 <= s1008;
      s1010 <= s1009;
      s1011 <= s1010;
      s1012 <= s1011;
      s1013 <= s1012;
      s1014 <= s1013;
      s1015 <= s1014;
      s1016 <= s1015;
      s1017 <= s1016;
      s1018 <= s1017;
      s1019 <= s1018;
      s1020 <= s1019;
      s1021 <= s1020;
      s1022 <= s1021;
      s1023 <= s1022;
      s1024 <= s1023;
      s1025 <= s1024;
      s1026 <= s1025;
      s1027 <= s1026;
      s1028 <= s1027;
      s1029 <= s1028;
      s1030 <= s1029;
      s1031 <= s1030;
      s1032 <= s1031;
      s1033 <= s1032;
      s1034 <= s1033;
      s1035 <= s1034;
      s1036 <= s1035;
      s1037 <= s1036;
      s1038 <= s1037;
      s1039 <= s1038;
      s1040 <= s1039;
      s1041 <= s1040;
      s1042 <= s1041;
      s1043 <= s1042;
      s1044 <= s1043;
      s1045 <= s1044;
      s1046 <= s1045;
      s1047 <= s1046;
      s1048 <= s1047;
      s1049 <= s1048;
      s1050 <= s1049;
      s1051 <= s1050;
      s1052 <= s1051;
      s1053 <= s1052;
      s1054 <= s1053;
      s1055 <= s1054;
      s1056 <= s1055;
      s1057 <= s1056;
      s1058 <= s1057;
      s1059 <= s1058;
      s1060 <= s1059;
      s1061 <= s1060;
      s1062 <= s1061;
      s1063 <= s1062;
      s1064 <= s1063;
      s1065 <= s1064;
      s1066 <= s1065;
      s1067 <= s1066;
      s1068 <= s1067;
      s1069 <= s1068;
      s1070 <= s1069;
      s1071 <= s1070;
      s1072 <= s1071;
      s1073 <= s1072;
      s1074 <= s1073;
      s1075 <= s1074;
      s1076 <= s1075;
      s1077 <= s1076;
      s1078 <= s1077;
      s1079 <= s1078;
      s1080 <= s1079;
      Y <= s1080;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_162_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 162 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_162_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_162_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      Y <= s161;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_246_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 246 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_246_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_246_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      Y <= s245;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_296_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 296 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_296_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_296_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      Y <= s295;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_365_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 365 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_365_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_365_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      Y <= s364;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_439_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 439 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_439_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_439_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      Y <= s438;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_507_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 507 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_507_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_507_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      Y <= s506;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_558_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 558 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_558_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_558_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      Y <= s557;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_624_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 624 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_624_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_624_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
signal s558 : std_logic_vector(33 downto 0) := (others => '0');
signal s559 : std_logic_vector(33 downto 0) := (others => '0');
signal s560 : std_logic_vector(33 downto 0) := (others => '0');
signal s561 : std_logic_vector(33 downto 0) := (others => '0');
signal s562 : std_logic_vector(33 downto 0) := (others => '0');
signal s563 : std_logic_vector(33 downto 0) := (others => '0');
signal s564 : std_logic_vector(33 downto 0) := (others => '0');
signal s565 : std_logic_vector(33 downto 0) := (others => '0');
signal s566 : std_logic_vector(33 downto 0) := (others => '0');
signal s567 : std_logic_vector(33 downto 0) := (others => '0');
signal s568 : std_logic_vector(33 downto 0) := (others => '0');
signal s569 : std_logic_vector(33 downto 0) := (others => '0');
signal s570 : std_logic_vector(33 downto 0) := (others => '0');
signal s571 : std_logic_vector(33 downto 0) := (others => '0');
signal s572 : std_logic_vector(33 downto 0) := (others => '0');
signal s573 : std_logic_vector(33 downto 0) := (others => '0');
signal s574 : std_logic_vector(33 downto 0) := (others => '0');
signal s575 : std_logic_vector(33 downto 0) := (others => '0');
signal s576 : std_logic_vector(33 downto 0) := (others => '0');
signal s577 : std_logic_vector(33 downto 0) := (others => '0');
signal s578 : std_logic_vector(33 downto 0) := (others => '0');
signal s579 : std_logic_vector(33 downto 0) := (others => '0');
signal s580 : std_logic_vector(33 downto 0) := (others => '0');
signal s581 : std_logic_vector(33 downto 0) := (others => '0');
signal s582 : std_logic_vector(33 downto 0) := (others => '0');
signal s583 : std_logic_vector(33 downto 0) := (others => '0');
signal s584 : std_logic_vector(33 downto 0) := (others => '0');
signal s585 : std_logic_vector(33 downto 0) := (others => '0');
signal s586 : std_logic_vector(33 downto 0) := (others => '0');
signal s587 : std_logic_vector(33 downto 0) := (others => '0');
signal s588 : std_logic_vector(33 downto 0) := (others => '0');
signal s589 : std_logic_vector(33 downto 0) := (others => '0');
signal s590 : std_logic_vector(33 downto 0) := (others => '0');
signal s591 : std_logic_vector(33 downto 0) := (others => '0');
signal s592 : std_logic_vector(33 downto 0) := (others => '0');
signal s593 : std_logic_vector(33 downto 0) := (others => '0');
signal s594 : std_logic_vector(33 downto 0) := (others => '0');
signal s595 : std_logic_vector(33 downto 0) := (others => '0');
signal s596 : std_logic_vector(33 downto 0) := (others => '0');
signal s597 : std_logic_vector(33 downto 0) := (others => '0');
signal s598 : std_logic_vector(33 downto 0) := (others => '0');
signal s599 : std_logic_vector(33 downto 0) := (others => '0');
signal s600 : std_logic_vector(33 downto 0) := (others => '0');
signal s601 : std_logic_vector(33 downto 0) := (others => '0');
signal s602 : std_logic_vector(33 downto 0) := (others => '0');
signal s603 : std_logic_vector(33 downto 0) := (others => '0');
signal s604 : std_logic_vector(33 downto 0) := (others => '0');
signal s605 : std_logic_vector(33 downto 0) := (others => '0');
signal s606 : std_logic_vector(33 downto 0) := (others => '0');
signal s607 : std_logic_vector(33 downto 0) := (others => '0');
signal s608 : std_logic_vector(33 downto 0) := (others => '0');
signal s609 : std_logic_vector(33 downto 0) := (others => '0');
signal s610 : std_logic_vector(33 downto 0) := (others => '0');
signal s611 : std_logic_vector(33 downto 0) := (others => '0');
signal s612 : std_logic_vector(33 downto 0) := (others => '0');
signal s613 : std_logic_vector(33 downto 0) := (others => '0');
signal s614 : std_logic_vector(33 downto 0) := (others => '0');
signal s615 : std_logic_vector(33 downto 0) := (others => '0');
signal s616 : std_logic_vector(33 downto 0) := (others => '0');
signal s617 : std_logic_vector(33 downto 0) := (others => '0');
signal s618 : std_logic_vector(33 downto 0) := (others => '0');
signal s619 : std_logic_vector(33 downto 0) := (others => '0');
signal s620 : std_logic_vector(33 downto 0) := (others => '0');
signal s621 : std_logic_vector(33 downto 0) := (others => '0');
signal s622 : std_logic_vector(33 downto 0) := (others => '0');
signal s623 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
      s558 <= "0000000000000000000000000000000000";
      s559 <= "0000000000000000000000000000000000";
      s560 <= "0000000000000000000000000000000000";
      s561 <= "0000000000000000000000000000000000";
      s562 <= "0000000000000000000000000000000000";
      s563 <= "0000000000000000000000000000000000";
      s564 <= "0000000000000000000000000000000000";
      s565 <= "0000000000000000000000000000000000";
      s566 <= "0000000000000000000000000000000000";
      s567 <= "0000000000000000000000000000000000";
      s568 <= "0000000000000000000000000000000000";
      s569 <= "0000000000000000000000000000000000";
      s570 <= "0000000000000000000000000000000000";
      s571 <= "0000000000000000000000000000000000";
      s572 <= "0000000000000000000000000000000000";
      s573 <= "0000000000000000000000000000000000";
      s574 <= "0000000000000000000000000000000000";
      s575 <= "0000000000000000000000000000000000";
      s576 <= "0000000000000000000000000000000000";
      s577 <= "0000000000000000000000000000000000";
      s578 <= "0000000000000000000000000000000000";
      s579 <= "0000000000000000000000000000000000";
      s580 <= "0000000000000000000000000000000000";
      s581 <= "0000000000000000000000000000000000";
      s582 <= "0000000000000000000000000000000000";
      s583 <= "0000000000000000000000000000000000";
      s584 <= "0000000000000000000000000000000000";
      s585 <= "0000000000000000000000000000000000";
      s586 <= "0000000000000000000000000000000000";
      s587 <= "0000000000000000000000000000000000";
      s588 <= "0000000000000000000000000000000000";
      s589 <= "0000000000000000000000000000000000";
      s590 <= "0000000000000000000000000000000000";
      s591 <= "0000000000000000000000000000000000";
      s592 <= "0000000000000000000000000000000000";
      s593 <= "0000000000000000000000000000000000";
      s594 <= "0000000000000000000000000000000000";
      s595 <= "0000000000000000000000000000000000";
      s596 <= "0000000000000000000000000000000000";
      s597 <= "0000000000000000000000000000000000";
      s598 <= "0000000000000000000000000000000000";
      s599 <= "0000000000000000000000000000000000";
      s600 <= "0000000000000000000000000000000000";
      s601 <= "0000000000000000000000000000000000";
      s602 <= "0000000000000000000000000000000000";
      s603 <= "0000000000000000000000000000000000";
      s604 <= "0000000000000000000000000000000000";
      s605 <= "0000000000000000000000000000000000";
      s606 <= "0000000000000000000000000000000000";
      s607 <= "0000000000000000000000000000000000";
      s608 <= "0000000000000000000000000000000000";
      s609 <= "0000000000000000000000000000000000";
      s610 <= "0000000000000000000000000000000000";
      s611 <= "0000000000000000000000000000000000";
      s612 <= "0000000000000000000000000000000000";
      s613 <= "0000000000000000000000000000000000";
      s614 <= "0000000000000000000000000000000000";
      s615 <= "0000000000000000000000000000000000";
      s616 <= "0000000000000000000000000000000000";
      s617 <= "0000000000000000000000000000000000";
      s618 <= "0000000000000000000000000000000000";
      s619 <= "0000000000000000000000000000000000";
      s620 <= "0000000000000000000000000000000000";
      s621 <= "0000000000000000000000000000000000";
      s622 <= "0000000000000000000000000000000000";
      s623 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      s558 <= s557;
      s559 <= s558;
      s560 <= s559;
      s561 <= s560;
      s562 <= s561;
      s563 <= s562;
      s564 <= s563;
      s565 <= s564;
      s566 <= s565;
      s567 <= s566;
      s568 <= s567;
      s569 <= s568;
      s570 <= s569;
      s571 <= s570;
      s572 <= s571;
      s573 <= s572;
      s574 <= s573;
      s575 <= s574;
      s576 <= s575;
      s577 <= s576;
      s578 <= s577;
      s579 <= s578;
      s580 <= s579;
      s581 <= s580;
      s582 <= s581;
      s583 <= s582;
      s584 <= s583;
      s585 <= s584;
      s586 <= s585;
      s587 <= s586;
      s588 <= s587;
      s589 <= s588;
      s590 <= s589;
      s591 <= s590;
      s592 <= s591;
      s593 <= s592;
      s594 <= s593;
      s595 <= s594;
      s596 <= s595;
      s597 <= s596;
      s598 <= s597;
      s599 <= s598;
      s600 <= s599;
      s601 <= s600;
      s602 <= s601;
      s603 <= s602;
      s604 <= s603;
      s605 <= s604;
      s606 <= s605;
      s607 <= s606;
      s608 <= s607;
      s609 <= s608;
      s610 <= s609;
      s611 <= s610;
      s612 <= s611;
      s613 <= s612;
      s614 <= s613;
      s615 <= s614;
      s616 <= s615;
      s617 <= s616;
      s618 <= s617;
      s619 <= s618;
      s620 <= s619;
      s621 <= s620;
      s622 <= s621;
      s623 <= s622;
      Y <= s623;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_73_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 73 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_73_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_73_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      Y <= s72;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 66 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      Y <= s65;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_75_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 75 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_75_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_75_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      Y <= s74;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 55 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      Y <= s54;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_70_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 70 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_70_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_70_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      Y <= s69;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 65 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      Y <= s64;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 67 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      Y <= s66;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_130_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 130 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_130_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_130_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      Y <= s129;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 97 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      Y <= s96;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_681_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 681 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_681_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_681_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
signal s558 : std_logic_vector(33 downto 0) := (others => '0');
signal s559 : std_logic_vector(33 downto 0) := (others => '0');
signal s560 : std_logic_vector(33 downto 0) := (others => '0');
signal s561 : std_logic_vector(33 downto 0) := (others => '0');
signal s562 : std_logic_vector(33 downto 0) := (others => '0');
signal s563 : std_logic_vector(33 downto 0) := (others => '0');
signal s564 : std_logic_vector(33 downto 0) := (others => '0');
signal s565 : std_logic_vector(33 downto 0) := (others => '0');
signal s566 : std_logic_vector(33 downto 0) := (others => '0');
signal s567 : std_logic_vector(33 downto 0) := (others => '0');
signal s568 : std_logic_vector(33 downto 0) := (others => '0');
signal s569 : std_logic_vector(33 downto 0) := (others => '0');
signal s570 : std_logic_vector(33 downto 0) := (others => '0');
signal s571 : std_logic_vector(33 downto 0) := (others => '0');
signal s572 : std_logic_vector(33 downto 0) := (others => '0');
signal s573 : std_logic_vector(33 downto 0) := (others => '0');
signal s574 : std_logic_vector(33 downto 0) := (others => '0');
signal s575 : std_logic_vector(33 downto 0) := (others => '0');
signal s576 : std_logic_vector(33 downto 0) := (others => '0');
signal s577 : std_logic_vector(33 downto 0) := (others => '0');
signal s578 : std_logic_vector(33 downto 0) := (others => '0');
signal s579 : std_logic_vector(33 downto 0) := (others => '0');
signal s580 : std_logic_vector(33 downto 0) := (others => '0');
signal s581 : std_logic_vector(33 downto 0) := (others => '0');
signal s582 : std_logic_vector(33 downto 0) := (others => '0');
signal s583 : std_logic_vector(33 downto 0) := (others => '0');
signal s584 : std_logic_vector(33 downto 0) := (others => '0');
signal s585 : std_logic_vector(33 downto 0) := (others => '0');
signal s586 : std_logic_vector(33 downto 0) := (others => '0');
signal s587 : std_logic_vector(33 downto 0) := (others => '0');
signal s588 : std_logic_vector(33 downto 0) := (others => '0');
signal s589 : std_logic_vector(33 downto 0) := (others => '0');
signal s590 : std_logic_vector(33 downto 0) := (others => '0');
signal s591 : std_logic_vector(33 downto 0) := (others => '0');
signal s592 : std_logic_vector(33 downto 0) := (others => '0');
signal s593 : std_logic_vector(33 downto 0) := (others => '0');
signal s594 : std_logic_vector(33 downto 0) := (others => '0');
signal s595 : std_logic_vector(33 downto 0) := (others => '0');
signal s596 : std_logic_vector(33 downto 0) := (others => '0');
signal s597 : std_logic_vector(33 downto 0) := (others => '0');
signal s598 : std_logic_vector(33 downto 0) := (others => '0');
signal s599 : std_logic_vector(33 downto 0) := (others => '0');
signal s600 : std_logic_vector(33 downto 0) := (others => '0');
signal s601 : std_logic_vector(33 downto 0) := (others => '0');
signal s602 : std_logic_vector(33 downto 0) := (others => '0');
signal s603 : std_logic_vector(33 downto 0) := (others => '0');
signal s604 : std_logic_vector(33 downto 0) := (others => '0');
signal s605 : std_logic_vector(33 downto 0) := (others => '0');
signal s606 : std_logic_vector(33 downto 0) := (others => '0');
signal s607 : std_logic_vector(33 downto 0) := (others => '0');
signal s608 : std_logic_vector(33 downto 0) := (others => '0');
signal s609 : std_logic_vector(33 downto 0) := (others => '0');
signal s610 : std_logic_vector(33 downto 0) := (others => '0');
signal s611 : std_logic_vector(33 downto 0) := (others => '0');
signal s612 : std_logic_vector(33 downto 0) := (others => '0');
signal s613 : std_logic_vector(33 downto 0) := (others => '0');
signal s614 : std_logic_vector(33 downto 0) := (others => '0');
signal s615 : std_logic_vector(33 downto 0) := (others => '0');
signal s616 : std_logic_vector(33 downto 0) := (others => '0');
signal s617 : std_logic_vector(33 downto 0) := (others => '0');
signal s618 : std_logic_vector(33 downto 0) := (others => '0');
signal s619 : std_logic_vector(33 downto 0) := (others => '0');
signal s620 : std_logic_vector(33 downto 0) := (others => '0');
signal s621 : std_logic_vector(33 downto 0) := (others => '0');
signal s622 : std_logic_vector(33 downto 0) := (others => '0');
signal s623 : std_logic_vector(33 downto 0) := (others => '0');
signal s624 : std_logic_vector(33 downto 0) := (others => '0');
signal s625 : std_logic_vector(33 downto 0) := (others => '0');
signal s626 : std_logic_vector(33 downto 0) := (others => '0');
signal s627 : std_logic_vector(33 downto 0) := (others => '0');
signal s628 : std_logic_vector(33 downto 0) := (others => '0');
signal s629 : std_logic_vector(33 downto 0) := (others => '0');
signal s630 : std_logic_vector(33 downto 0) := (others => '0');
signal s631 : std_logic_vector(33 downto 0) := (others => '0');
signal s632 : std_logic_vector(33 downto 0) := (others => '0');
signal s633 : std_logic_vector(33 downto 0) := (others => '0');
signal s634 : std_logic_vector(33 downto 0) := (others => '0');
signal s635 : std_logic_vector(33 downto 0) := (others => '0');
signal s636 : std_logic_vector(33 downto 0) := (others => '0');
signal s637 : std_logic_vector(33 downto 0) := (others => '0');
signal s638 : std_logic_vector(33 downto 0) := (others => '0');
signal s639 : std_logic_vector(33 downto 0) := (others => '0');
signal s640 : std_logic_vector(33 downto 0) := (others => '0');
signal s641 : std_logic_vector(33 downto 0) := (others => '0');
signal s642 : std_logic_vector(33 downto 0) := (others => '0');
signal s643 : std_logic_vector(33 downto 0) := (others => '0');
signal s644 : std_logic_vector(33 downto 0) := (others => '0');
signal s645 : std_logic_vector(33 downto 0) := (others => '0');
signal s646 : std_logic_vector(33 downto 0) := (others => '0');
signal s647 : std_logic_vector(33 downto 0) := (others => '0');
signal s648 : std_logic_vector(33 downto 0) := (others => '0');
signal s649 : std_logic_vector(33 downto 0) := (others => '0');
signal s650 : std_logic_vector(33 downto 0) := (others => '0');
signal s651 : std_logic_vector(33 downto 0) := (others => '0');
signal s652 : std_logic_vector(33 downto 0) := (others => '0');
signal s653 : std_logic_vector(33 downto 0) := (others => '0');
signal s654 : std_logic_vector(33 downto 0) := (others => '0');
signal s655 : std_logic_vector(33 downto 0) := (others => '0');
signal s656 : std_logic_vector(33 downto 0) := (others => '0');
signal s657 : std_logic_vector(33 downto 0) := (others => '0');
signal s658 : std_logic_vector(33 downto 0) := (others => '0');
signal s659 : std_logic_vector(33 downto 0) := (others => '0');
signal s660 : std_logic_vector(33 downto 0) := (others => '0');
signal s661 : std_logic_vector(33 downto 0) := (others => '0');
signal s662 : std_logic_vector(33 downto 0) := (others => '0');
signal s663 : std_logic_vector(33 downto 0) := (others => '0');
signal s664 : std_logic_vector(33 downto 0) := (others => '0');
signal s665 : std_logic_vector(33 downto 0) := (others => '0');
signal s666 : std_logic_vector(33 downto 0) := (others => '0');
signal s667 : std_logic_vector(33 downto 0) := (others => '0');
signal s668 : std_logic_vector(33 downto 0) := (others => '0');
signal s669 : std_logic_vector(33 downto 0) := (others => '0');
signal s670 : std_logic_vector(33 downto 0) := (others => '0');
signal s671 : std_logic_vector(33 downto 0) := (others => '0');
signal s672 : std_logic_vector(33 downto 0) := (others => '0');
signal s673 : std_logic_vector(33 downto 0) := (others => '0');
signal s674 : std_logic_vector(33 downto 0) := (others => '0');
signal s675 : std_logic_vector(33 downto 0) := (others => '0');
signal s676 : std_logic_vector(33 downto 0) := (others => '0');
signal s677 : std_logic_vector(33 downto 0) := (others => '0');
signal s678 : std_logic_vector(33 downto 0) := (others => '0');
signal s679 : std_logic_vector(33 downto 0) := (others => '0');
signal s680 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
      s558 <= "0000000000000000000000000000000000";
      s559 <= "0000000000000000000000000000000000";
      s560 <= "0000000000000000000000000000000000";
      s561 <= "0000000000000000000000000000000000";
      s562 <= "0000000000000000000000000000000000";
      s563 <= "0000000000000000000000000000000000";
      s564 <= "0000000000000000000000000000000000";
      s565 <= "0000000000000000000000000000000000";
      s566 <= "0000000000000000000000000000000000";
      s567 <= "0000000000000000000000000000000000";
      s568 <= "0000000000000000000000000000000000";
      s569 <= "0000000000000000000000000000000000";
      s570 <= "0000000000000000000000000000000000";
      s571 <= "0000000000000000000000000000000000";
      s572 <= "0000000000000000000000000000000000";
      s573 <= "0000000000000000000000000000000000";
      s574 <= "0000000000000000000000000000000000";
      s575 <= "0000000000000000000000000000000000";
      s576 <= "0000000000000000000000000000000000";
      s577 <= "0000000000000000000000000000000000";
      s578 <= "0000000000000000000000000000000000";
      s579 <= "0000000000000000000000000000000000";
      s580 <= "0000000000000000000000000000000000";
      s581 <= "0000000000000000000000000000000000";
      s582 <= "0000000000000000000000000000000000";
      s583 <= "0000000000000000000000000000000000";
      s584 <= "0000000000000000000000000000000000";
      s585 <= "0000000000000000000000000000000000";
      s586 <= "0000000000000000000000000000000000";
      s587 <= "0000000000000000000000000000000000";
      s588 <= "0000000000000000000000000000000000";
      s589 <= "0000000000000000000000000000000000";
      s590 <= "0000000000000000000000000000000000";
      s591 <= "0000000000000000000000000000000000";
      s592 <= "0000000000000000000000000000000000";
      s593 <= "0000000000000000000000000000000000";
      s594 <= "0000000000000000000000000000000000";
      s595 <= "0000000000000000000000000000000000";
      s596 <= "0000000000000000000000000000000000";
      s597 <= "0000000000000000000000000000000000";
      s598 <= "0000000000000000000000000000000000";
      s599 <= "0000000000000000000000000000000000";
      s600 <= "0000000000000000000000000000000000";
      s601 <= "0000000000000000000000000000000000";
      s602 <= "0000000000000000000000000000000000";
      s603 <= "0000000000000000000000000000000000";
      s604 <= "0000000000000000000000000000000000";
      s605 <= "0000000000000000000000000000000000";
      s606 <= "0000000000000000000000000000000000";
      s607 <= "0000000000000000000000000000000000";
      s608 <= "0000000000000000000000000000000000";
      s609 <= "0000000000000000000000000000000000";
      s610 <= "0000000000000000000000000000000000";
      s611 <= "0000000000000000000000000000000000";
      s612 <= "0000000000000000000000000000000000";
      s613 <= "0000000000000000000000000000000000";
      s614 <= "0000000000000000000000000000000000";
      s615 <= "0000000000000000000000000000000000";
      s616 <= "0000000000000000000000000000000000";
      s617 <= "0000000000000000000000000000000000";
      s618 <= "0000000000000000000000000000000000";
      s619 <= "0000000000000000000000000000000000";
      s620 <= "0000000000000000000000000000000000";
      s621 <= "0000000000000000000000000000000000";
      s622 <= "0000000000000000000000000000000000";
      s623 <= "0000000000000000000000000000000000";
      s624 <= "0000000000000000000000000000000000";
      s625 <= "0000000000000000000000000000000000";
      s626 <= "0000000000000000000000000000000000";
      s627 <= "0000000000000000000000000000000000";
      s628 <= "0000000000000000000000000000000000";
      s629 <= "0000000000000000000000000000000000";
      s630 <= "0000000000000000000000000000000000";
      s631 <= "0000000000000000000000000000000000";
      s632 <= "0000000000000000000000000000000000";
      s633 <= "0000000000000000000000000000000000";
      s634 <= "0000000000000000000000000000000000";
      s635 <= "0000000000000000000000000000000000";
      s636 <= "0000000000000000000000000000000000";
      s637 <= "0000000000000000000000000000000000";
      s638 <= "0000000000000000000000000000000000";
      s639 <= "0000000000000000000000000000000000";
      s640 <= "0000000000000000000000000000000000";
      s641 <= "0000000000000000000000000000000000";
      s642 <= "0000000000000000000000000000000000";
      s643 <= "0000000000000000000000000000000000";
      s644 <= "0000000000000000000000000000000000";
      s645 <= "0000000000000000000000000000000000";
      s646 <= "0000000000000000000000000000000000";
      s647 <= "0000000000000000000000000000000000";
      s648 <= "0000000000000000000000000000000000";
      s649 <= "0000000000000000000000000000000000";
      s650 <= "0000000000000000000000000000000000";
      s651 <= "0000000000000000000000000000000000";
      s652 <= "0000000000000000000000000000000000";
      s653 <= "0000000000000000000000000000000000";
      s654 <= "0000000000000000000000000000000000";
      s655 <= "0000000000000000000000000000000000";
      s656 <= "0000000000000000000000000000000000";
      s657 <= "0000000000000000000000000000000000";
      s658 <= "0000000000000000000000000000000000";
      s659 <= "0000000000000000000000000000000000";
      s660 <= "0000000000000000000000000000000000";
      s661 <= "0000000000000000000000000000000000";
      s662 <= "0000000000000000000000000000000000";
      s663 <= "0000000000000000000000000000000000";
      s664 <= "0000000000000000000000000000000000";
      s665 <= "0000000000000000000000000000000000";
      s666 <= "0000000000000000000000000000000000";
      s667 <= "0000000000000000000000000000000000";
      s668 <= "0000000000000000000000000000000000";
      s669 <= "0000000000000000000000000000000000";
      s670 <= "0000000000000000000000000000000000";
      s671 <= "0000000000000000000000000000000000";
      s672 <= "0000000000000000000000000000000000";
      s673 <= "0000000000000000000000000000000000";
      s674 <= "0000000000000000000000000000000000";
      s675 <= "0000000000000000000000000000000000";
      s676 <= "0000000000000000000000000000000000";
      s677 <= "0000000000000000000000000000000000";
      s678 <= "0000000000000000000000000000000000";
      s679 <= "0000000000000000000000000000000000";
      s680 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      s558 <= s557;
      s559 <= s558;
      s560 <= s559;
      s561 <= s560;
      s562 <= s561;
      s563 <= s562;
      s564 <= s563;
      s565 <= s564;
      s566 <= s565;
      s567 <= s566;
      s568 <= s567;
      s569 <= s568;
      s570 <= s569;
      s571 <= s570;
      s572 <= s571;
      s573 <= s572;
      s574 <= s573;
      s575 <= s574;
      s576 <= s575;
      s577 <= s576;
      s578 <= s577;
      s579 <= s578;
      s580 <= s579;
      s581 <= s580;
      s582 <= s581;
      s583 <= s582;
      s584 <= s583;
      s585 <= s584;
      s586 <= s585;
      s587 <= s586;
      s588 <= s587;
      s589 <= s588;
      s590 <= s589;
      s591 <= s590;
      s592 <= s591;
      s593 <= s592;
      s594 <= s593;
      s595 <= s594;
      s596 <= s595;
      s597 <= s596;
      s598 <= s597;
      s599 <= s598;
      s600 <= s599;
      s601 <= s600;
      s602 <= s601;
      s603 <= s602;
      s604 <= s603;
      s605 <= s604;
      s606 <= s605;
      s607 <= s606;
      s608 <= s607;
      s609 <= s608;
      s610 <= s609;
      s611 <= s610;
      s612 <= s611;
      s613 <= s612;
      s614 <= s613;
      s615 <= s614;
      s616 <= s615;
      s617 <= s616;
      s618 <= s617;
      s619 <= s618;
      s620 <= s619;
      s621 <= s620;
      s622 <= s621;
      s623 <= s622;
      s624 <= s623;
      s625 <= s624;
      s626 <= s625;
      s627 <= s626;
      s628 <= s627;
      s629 <= s628;
      s630 <= s629;
      s631 <= s630;
      s632 <= s631;
      s633 <= s632;
      s634 <= s633;
      s635 <= s634;
      s636 <= s635;
      s637 <= s636;
      s638 <= s637;
      s639 <= s638;
      s640 <= s639;
      s641 <= s640;
      s642 <= s641;
      s643 <= s642;
      s644 <= s643;
      s645 <= s644;
      s646 <= s645;
      s647 <= s646;
      s648 <= s647;
      s649 <= s648;
      s650 <= s649;
      s651 <= s650;
      s652 <= s651;
      s653 <= s652;
      s654 <= s653;
      s655 <= s654;
      s656 <= s655;
      s657 <= s656;
      s658 <= s657;
      s659 <= s658;
      s660 <= s659;
      s661 <= s660;
      s662 <= s661;
      s663 <= s662;
      s664 <= s663;
      s665 <= s664;
      s666 <= s665;
      s667 <= s666;
      s668 <= s667;
      s669 <= s668;
      s670 <= s669;
      s671 <= s670;
      s672 <= s671;
      s673 <= s672;
      s674 <= s673;
      s675 <= s674;
      s676 <= s675;
      s677 <= s676;
      s678 <= s677;
      s679 <= s678;
      s680 <= s679;
      Y <= s680;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_735_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 735 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_735_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_735_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
signal s558 : std_logic_vector(33 downto 0) := (others => '0');
signal s559 : std_logic_vector(33 downto 0) := (others => '0');
signal s560 : std_logic_vector(33 downto 0) := (others => '0');
signal s561 : std_logic_vector(33 downto 0) := (others => '0');
signal s562 : std_logic_vector(33 downto 0) := (others => '0');
signal s563 : std_logic_vector(33 downto 0) := (others => '0');
signal s564 : std_logic_vector(33 downto 0) := (others => '0');
signal s565 : std_logic_vector(33 downto 0) := (others => '0');
signal s566 : std_logic_vector(33 downto 0) := (others => '0');
signal s567 : std_logic_vector(33 downto 0) := (others => '0');
signal s568 : std_logic_vector(33 downto 0) := (others => '0');
signal s569 : std_logic_vector(33 downto 0) := (others => '0');
signal s570 : std_logic_vector(33 downto 0) := (others => '0');
signal s571 : std_logic_vector(33 downto 0) := (others => '0');
signal s572 : std_logic_vector(33 downto 0) := (others => '0');
signal s573 : std_logic_vector(33 downto 0) := (others => '0');
signal s574 : std_logic_vector(33 downto 0) := (others => '0');
signal s575 : std_logic_vector(33 downto 0) := (others => '0');
signal s576 : std_logic_vector(33 downto 0) := (others => '0');
signal s577 : std_logic_vector(33 downto 0) := (others => '0');
signal s578 : std_logic_vector(33 downto 0) := (others => '0');
signal s579 : std_logic_vector(33 downto 0) := (others => '0');
signal s580 : std_logic_vector(33 downto 0) := (others => '0');
signal s581 : std_logic_vector(33 downto 0) := (others => '0');
signal s582 : std_logic_vector(33 downto 0) := (others => '0');
signal s583 : std_logic_vector(33 downto 0) := (others => '0');
signal s584 : std_logic_vector(33 downto 0) := (others => '0');
signal s585 : std_logic_vector(33 downto 0) := (others => '0');
signal s586 : std_logic_vector(33 downto 0) := (others => '0');
signal s587 : std_logic_vector(33 downto 0) := (others => '0');
signal s588 : std_logic_vector(33 downto 0) := (others => '0');
signal s589 : std_logic_vector(33 downto 0) := (others => '0');
signal s590 : std_logic_vector(33 downto 0) := (others => '0');
signal s591 : std_logic_vector(33 downto 0) := (others => '0');
signal s592 : std_logic_vector(33 downto 0) := (others => '0');
signal s593 : std_logic_vector(33 downto 0) := (others => '0');
signal s594 : std_logic_vector(33 downto 0) := (others => '0');
signal s595 : std_logic_vector(33 downto 0) := (others => '0');
signal s596 : std_logic_vector(33 downto 0) := (others => '0');
signal s597 : std_logic_vector(33 downto 0) := (others => '0');
signal s598 : std_logic_vector(33 downto 0) := (others => '0');
signal s599 : std_logic_vector(33 downto 0) := (others => '0');
signal s600 : std_logic_vector(33 downto 0) := (others => '0');
signal s601 : std_logic_vector(33 downto 0) := (others => '0');
signal s602 : std_logic_vector(33 downto 0) := (others => '0');
signal s603 : std_logic_vector(33 downto 0) := (others => '0');
signal s604 : std_logic_vector(33 downto 0) := (others => '0');
signal s605 : std_logic_vector(33 downto 0) := (others => '0');
signal s606 : std_logic_vector(33 downto 0) := (others => '0');
signal s607 : std_logic_vector(33 downto 0) := (others => '0');
signal s608 : std_logic_vector(33 downto 0) := (others => '0');
signal s609 : std_logic_vector(33 downto 0) := (others => '0');
signal s610 : std_logic_vector(33 downto 0) := (others => '0');
signal s611 : std_logic_vector(33 downto 0) := (others => '0');
signal s612 : std_logic_vector(33 downto 0) := (others => '0');
signal s613 : std_logic_vector(33 downto 0) := (others => '0');
signal s614 : std_logic_vector(33 downto 0) := (others => '0');
signal s615 : std_logic_vector(33 downto 0) := (others => '0');
signal s616 : std_logic_vector(33 downto 0) := (others => '0');
signal s617 : std_logic_vector(33 downto 0) := (others => '0');
signal s618 : std_logic_vector(33 downto 0) := (others => '0');
signal s619 : std_logic_vector(33 downto 0) := (others => '0');
signal s620 : std_logic_vector(33 downto 0) := (others => '0');
signal s621 : std_logic_vector(33 downto 0) := (others => '0');
signal s622 : std_logic_vector(33 downto 0) := (others => '0');
signal s623 : std_logic_vector(33 downto 0) := (others => '0');
signal s624 : std_logic_vector(33 downto 0) := (others => '0');
signal s625 : std_logic_vector(33 downto 0) := (others => '0');
signal s626 : std_logic_vector(33 downto 0) := (others => '0');
signal s627 : std_logic_vector(33 downto 0) := (others => '0');
signal s628 : std_logic_vector(33 downto 0) := (others => '0');
signal s629 : std_logic_vector(33 downto 0) := (others => '0');
signal s630 : std_logic_vector(33 downto 0) := (others => '0');
signal s631 : std_logic_vector(33 downto 0) := (others => '0');
signal s632 : std_logic_vector(33 downto 0) := (others => '0');
signal s633 : std_logic_vector(33 downto 0) := (others => '0');
signal s634 : std_logic_vector(33 downto 0) := (others => '0');
signal s635 : std_logic_vector(33 downto 0) := (others => '0');
signal s636 : std_logic_vector(33 downto 0) := (others => '0');
signal s637 : std_logic_vector(33 downto 0) := (others => '0');
signal s638 : std_logic_vector(33 downto 0) := (others => '0');
signal s639 : std_logic_vector(33 downto 0) := (others => '0');
signal s640 : std_logic_vector(33 downto 0) := (others => '0');
signal s641 : std_logic_vector(33 downto 0) := (others => '0');
signal s642 : std_logic_vector(33 downto 0) := (others => '0');
signal s643 : std_logic_vector(33 downto 0) := (others => '0');
signal s644 : std_logic_vector(33 downto 0) := (others => '0');
signal s645 : std_logic_vector(33 downto 0) := (others => '0');
signal s646 : std_logic_vector(33 downto 0) := (others => '0');
signal s647 : std_logic_vector(33 downto 0) := (others => '0');
signal s648 : std_logic_vector(33 downto 0) := (others => '0');
signal s649 : std_logic_vector(33 downto 0) := (others => '0');
signal s650 : std_logic_vector(33 downto 0) := (others => '0');
signal s651 : std_logic_vector(33 downto 0) := (others => '0');
signal s652 : std_logic_vector(33 downto 0) := (others => '0');
signal s653 : std_logic_vector(33 downto 0) := (others => '0');
signal s654 : std_logic_vector(33 downto 0) := (others => '0');
signal s655 : std_logic_vector(33 downto 0) := (others => '0');
signal s656 : std_logic_vector(33 downto 0) := (others => '0');
signal s657 : std_logic_vector(33 downto 0) := (others => '0');
signal s658 : std_logic_vector(33 downto 0) := (others => '0');
signal s659 : std_logic_vector(33 downto 0) := (others => '0');
signal s660 : std_logic_vector(33 downto 0) := (others => '0');
signal s661 : std_logic_vector(33 downto 0) := (others => '0');
signal s662 : std_logic_vector(33 downto 0) := (others => '0');
signal s663 : std_logic_vector(33 downto 0) := (others => '0');
signal s664 : std_logic_vector(33 downto 0) := (others => '0');
signal s665 : std_logic_vector(33 downto 0) := (others => '0');
signal s666 : std_logic_vector(33 downto 0) := (others => '0');
signal s667 : std_logic_vector(33 downto 0) := (others => '0');
signal s668 : std_logic_vector(33 downto 0) := (others => '0');
signal s669 : std_logic_vector(33 downto 0) := (others => '0');
signal s670 : std_logic_vector(33 downto 0) := (others => '0');
signal s671 : std_logic_vector(33 downto 0) := (others => '0');
signal s672 : std_logic_vector(33 downto 0) := (others => '0');
signal s673 : std_logic_vector(33 downto 0) := (others => '0');
signal s674 : std_logic_vector(33 downto 0) := (others => '0');
signal s675 : std_logic_vector(33 downto 0) := (others => '0');
signal s676 : std_logic_vector(33 downto 0) := (others => '0');
signal s677 : std_logic_vector(33 downto 0) := (others => '0');
signal s678 : std_logic_vector(33 downto 0) := (others => '0');
signal s679 : std_logic_vector(33 downto 0) := (others => '0');
signal s680 : std_logic_vector(33 downto 0) := (others => '0');
signal s681 : std_logic_vector(33 downto 0) := (others => '0');
signal s682 : std_logic_vector(33 downto 0) := (others => '0');
signal s683 : std_logic_vector(33 downto 0) := (others => '0');
signal s684 : std_logic_vector(33 downto 0) := (others => '0');
signal s685 : std_logic_vector(33 downto 0) := (others => '0');
signal s686 : std_logic_vector(33 downto 0) := (others => '0');
signal s687 : std_logic_vector(33 downto 0) := (others => '0');
signal s688 : std_logic_vector(33 downto 0) := (others => '0');
signal s689 : std_logic_vector(33 downto 0) := (others => '0');
signal s690 : std_logic_vector(33 downto 0) := (others => '0');
signal s691 : std_logic_vector(33 downto 0) := (others => '0');
signal s692 : std_logic_vector(33 downto 0) := (others => '0');
signal s693 : std_logic_vector(33 downto 0) := (others => '0');
signal s694 : std_logic_vector(33 downto 0) := (others => '0');
signal s695 : std_logic_vector(33 downto 0) := (others => '0');
signal s696 : std_logic_vector(33 downto 0) := (others => '0');
signal s697 : std_logic_vector(33 downto 0) := (others => '0');
signal s698 : std_logic_vector(33 downto 0) := (others => '0');
signal s699 : std_logic_vector(33 downto 0) := (others => '0');
signal s700 : std_logic_vector(33 downto 0) := (others => '0');
signal s701 : std_logic_vector(33 downto 0) := (others => '0');
signal s702 : std_logic_vector(33 downto 0) := (others => '0');
signal s703 : std_logic_vector(33 downto 0) := (others => '0');
signal s704 : std_logic_vector(33 downto 0) := (others => '0');
signal s705 : std_logic_vector(33 downto 0) := (others => '0');
signal s706 : std_logic_vector(33 downto 0) := (others => '0');
signal s707 : std_logic_vector(33 downto 0) := (others => '0');
signal s708 : std_logic_vector(33 downto 0) := (others => '0');
signal s709 : std_logic_vector(33 downto 0) := (others => '0');
signal s710 : std_logic_vector(33 downto 0) := (others => '0');
signal s711 : std_logic_vector(33 downto 0) := (others => '0');
signal s712 : std_logic_vector(33 downto 0) := (others => '0');
signal s713 : std_logic_vector(33 downto 0) := (others => '0');
signal s714 : std_logic_vector(33 downto 0) := (others => '0');
signal s715 : std_logic_vector(33 downto 0) := (others => '0');
signal s716 : std_logic_vector(33 downto 0) := (others => '0');
signal s717 : std_logic_vector(33 downto 0) := (others => '0');
signal s718 : std_logic_vector(33 downto 0) := (others => '0');
signal s719 : std_logic_vector(33 downto 0) := (others => '0');
signal s720 : std_logic_vector(33 downto 0) := (others => '0');
signal s721 : std_logic_vector(33 downto 0) := (others => '0');
signal s722 : std_logic_vector(33 downto 0) := (others => '0');
signal s723 : std_logic_vector(33 downto 0) := (others => '0');
signal s724 : std_logic_vector(33 downto 0) := (others => '0');
signal s725 : std_logic_vector(33 downto 0) := (others => '0');
signal s726 : std_logic_vector(33 downto 0) := (others => '0');
signal s727 : std_logic_vector(33 downto 0) := (others => '0');
signal s728 : std_logic_vector(33 downto 0) := (others => '0');
signal s729 : std_logic_vector(33 downto 0) := (others => '0');
signal s730 : std_logic_vector(33 downto 0) := (others => '0');
signal s731 : std_logic_vector(33 downto 0) := (others => '0');
signal s732 : std_logic_vector(33 downto 0) := (others => '0');
signal s733 : std_logic_vector(33 downto 0) := (others => '0');
signal s734 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
      s558 <= "0000000000000000000000000000000000";
      s559 <= "0000000000000000000000000000000000";
      s560 <= "0000000000000000000000000000000000";
      s561 <= "0000000000000000000000000000000000";
      s562 <= "0000000000000000000000000000000000";
      s563 <= "0000000000000000000000000000000000";
      s564 <= "0000000000000000000000000000000000";
      s565 <= "0000000000000000000000000000000000";
      s566 <= "0000000000000000000000000000000000";
      s567 <= "0000000000000000000000000000000000";
      s568 <= "0000000000000000000000000000000000";
      s569 <= "0000000000000000000000000000000000";
      s570 <= "0000000000000000000000000000000000";
      s571 <= "0000000000000000000000000000000000";
      s572 <= "0000000000000000000000000000000000";
      s573 <= "0000000000000000000000000000000000";
      s574 <= "0000000000000000000000000000000000";
      s575 <= "0000000000000000000000000000000000";
      s576 <= "0000000000000000000000000000000000";
      s577 <= "0000000000000000000000000000000000";
      s578 <= "0000000000000000000000000000000000";
      s579 <= "0000000000000000000000000000000000";
      s580 <= "0000000000000000000000000000000000";
      s581 <= "0000000000000000000000000000000000";
      s582 <= "0000000000000000000000000000000000";
      s583 <= "0000000000000000000000000000000000";
      s584 <= "0000000000000000000000000000000000";
      s585 <= "0000000000000000000000000000000000";
      s586 <= "0000000000000000000000000000000000";
      s587 <= "0000000000000000000000000000000000";
      s588 <= "0000000000000000000000000000000000";
      s589 <= "0000000000000000000000000000000000";
      s590 <= "0000000000000000000000000000000000";
      s591 <= "0000000000000000000000000000000000";
      s592 <= "0000000000000000000000000000000000";
      s593 <= "0000000000000000000000000000000000";
      s594 <= "0000000000000000000000000000000000";
      s595 <= "0000000000000000000000000000000000";
      s596 <= "0000000000000000000000000000000000";
      s597 <= "0000000000000000000000000000000000";
      s598 <= "0000000000000000000000000000000000";
      s599 <= "0000000000000000000000000000000000";
      s600 <= "0000000000000000000000000000000000";
      s601 <= "0000000000000000000000000000000000";
      s602 <= "0000000000000000000000000000000000";
      s603 <= "0000000000000000000000000000000000";
      s604 <= "0000000000000000000000000000000000";
      s605 <= "0000000000000000000000000000000000";
      s606 <= "0000000000000000000000000000000000";
      s607 <= "0000000000000000000000000000000000";
      s608 <= "0000000000000000000000000000000000";
      s609 <= "0000000000000000000000000000000000";
      s610 <= "0000000000000000000000000000000000";
      s611 <= "0000000000000000000000000000000000";
      s612 <= "0000000000000000000000000000000000";
      s613 <= "0000000000000000000000000000000000";
      s614 <= "0000000000000000000000000000000000";
      s615 <= "0000000000000000000000000000000000";
      s616 <= "0000000000000000000000000000000000";
      s617 <= "0000000000000000000000000000000000";
      s618 <= "0000000000000000000000000000000000";
      s619 <= "0000000000000000000000000000000000";
      s620 <= "0000000000000000000000000000000000";
      s621 <= "0000000000000000000000000000000000";
      s622 <= "0000000000000000000000000000000000";
      s623 <= "0000000000000000000000000000000000";
      s624 <= "0000000000000000000000000000000000";
      s625 <= "0000000000000000000000000000000000";
      s626 <= "0000000000000000000000000000000000";
      s627 <= "0000000000000000000000000000000000";
      s628 <= "0000000000000000000000000000000000";
      s629 <= "0000000000000000000000000000000000";
      s630 <= "0000000000000000000000000000000000";
      s631 <= "0000000000000000000000000000000000";
      s632 <= "0000000000000000000000000000000000";
      s633 <= "0000000000000000000000000000000000";
      s634 <= "0000000000000000000000000000000000";
      s635 <= "0000000000000000000000000000000000";
      s636 <= "0000000000000000000000000000000000";
      s637 <= "0000000000000000000000000000000000";
      s638 <= "0000000000000000000000000000000000";
      s639 <= "0000000000000000000000000000000000";
      s640 <= "0000000000000000000000000000000000";
      s641 <= "0000000000000000000000000000000000";
      s642 <= "0000000000000000000000000000000000";
      s643 <= "0000000000000000000000000000000000";
      s644 <= "0000000000000000000000000000000000";
      s645 <= "0000000000000000000000000000000000";
      s646 <= "0000000000000000000000000000000000";
      s647 <= "0000000000000000000000000000000000";
      s648 <= "0000000000000000000000000000000000";
      s649 <= "0000000000000000000000000000000000";
      s650 <= "0000000000000000000000000000000000";
      s651 <= "0000000000000000000000000000000000";
      s652 <= "0000000000000000000000000000000000";
      s653 <= "0000000000000000000000000000000000";
      s654 <= "0000000000000000000000000000000000";
      s655 <= "0000000000000000000000000000000000";
      s656 <= "0000000000000000000000000000000000";
      s657 <= "0000000000000000000000000000000000";
      s658 <= "0000000000000000000000000000000000";
      s659 <= "0000000000000000000000000000000000";
      s660 <= "0000000000000000000000000000000000";
      s661 <= "0000000000000000000000000000000000";
      s662 <= "0000000000000000000000000000000000";
      s663 <= "0000000000000000000000000000000000";
      s664 <= "0000000000000000000000000000000000";
      s665 <= "0000000000000000000000000000000000";
      s666 <= "0000000000000000000000000000000000";
      s667 <= "0000000000000000000000000000000000";
      s668 <= "0000000000000000000000000000000000";
      s669 <= "0000000000000000000000000000000000";
      s670 <= "0000000000000000000000000000000000";
      s671 <= "0000000000000000000000000000000000";
      s672 <= "0000000000000000000000000000000000";
      s673 <= "0000000000000000000000000000000000";
      s674 <= "0000000000000000000000000000000000";
      s675 <= "0000000000000000000000000000000000";
      s676 <= "0000000000000000000000000000000000";
      s677 <= "0000000000000000000000000000000000";
      s678 <= "0000000000000000000000000000000000";
      s679 <= "0000000000000000000000000000000000";
      s680 <= "0000000000000000000000000000000000";
      s681 <= "0000000000000000000000000000000000";
      s682 <= "0000000000000000000000000000000000";
      s683 <= "0000000000000000000000000000000000";
      s684 <= "0000000000000000000000000000000000";
      s685 <= "0000000000000000000000000000000000";
      s686 <= "0000000000000000000000000000000000";
      s687 <= "0000000000000000000000000000000000";
      s688 <= "0000000000000000000000000000000000";
      s689 <= "0000000000000000000000000000000000";
      s690 <= "0000000000000000000000000000000000";
      s691 <= "0000000000000000000000000000000000";
      s692 <= "0000000000000000000000000000000000";
      s693 <= "0000000000000000000000000000000000";
      s694 <= "0000000000000000000000000000000000";
      s695 <= "0000000000000000000000000000000000";
      s696 <= "0000000000000000000000000000000000";
      s697 <= "0000000000000000000000000000000000";
      s698 <= "0000000000000000000000000000000000";
      s699 <= "0000000000000000000000000000000000";
      s700 <= "0000000000000000000000000000000000";
      s701 <= "0000000000000000000000000000000000";
      s702 <= "0000000000000000000000000000000000";
      s703 <= "0000000000000000000000000000000000";
      s704 <= "0000000000000000000000000000000000";
      s705 <= "0000000000000000000000000000000000";
      s706 <= "0000000000000000000000000000000000";
      s707 <= "0000000000000000000000000000000000";
      s708 <= "0000000000000000000000000000000000";
      s709 <= "0000000000000000000000000000000000";
      s710 <= "0000000000000000000000000000000000";
      s711 <= "0000000000000000000000000000000000";
      s712 <= "0000000000000000000000000000000000";
      s713 <= "0000000000000000000000000000000000";
      s714 <= "0000000000000000000000000000000000";
      s715 <= "0000000000000000000000000000000000";
      s716 <= "0000000000000000000000000000000000";
      s717 <= "0000000000000000000000000000000000";
      s718 <= "0000000000000000000000000000000000";
      s719 <= "0000000000000000000000000000000000";
      s720 <= "0000000000000000000000000000000000";
      s721 <= "0000000000000000000000000000000000";
      s722 <= "0000000000000000000000000000000000";
      s723 <= "0000000000000000000000000000000000";
      s724 <= "0000000000000000000000000000000000";
      s725 <= "0000000000000000000000000000000000";
      s726 <= "0000000000000000000000000000000000";
      s727 <= "0000000000000000000000000000000000";
      s728 <= "0000000000000000000000000000000000";
      s729 <= "0000000000000000000000000000000000";
      s730 <= "0000000000000000000000000000000000";
      s731 <= "0000000000000000000000000000000000";
      s732 <= "0000000000000000000000000000000000";
      s733 <= "0000000000000000000000000000000000";
      s734 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      s558 <= s557;
      s559 <= s558;
      s560 <= s559;
      s561 <= s560;
      s562 <= s561;
      s563 <= s562;
      s564 <= s563;
      s565 <= s564;
      s566 <= s565;
      s567 <= s566;
      s568 <= s567;
      s569 <= s568;
      s570 <= s569;
      s571 <= s570;
      s572 <= s571;
      s573 <= s572;
      s574 <= s573;
      s575 <= s574;
      s576 <= s575;
      s577 <= s576;
      s578 <= s577;
      s579 <= s578;
      s580 <= s579;
      s581 <= s580;
      s582 <= s581;
      s583 <= s582;
      s584 <= s583;
      s585 <= s584;
      s586 <= s585;
      s587 <= s586;
      s588 <= s587;
      s589 <= s588;
      s590 <= s589;
      s591 <= s590;
      s592 <= s591;
      s593 <= s592;
      s594 <= s593;
      s595 <= s594;
      s596 <= s595;
      s597 <= s596;
      s598 <= s597;
      s599 <= s598;
      s600 <= s599;
      s601 <= s600;
      s602 <= s601;
      s603 <= s602;
      s604 <= s603;
      s605 <= s604;
      s606 <= s605;
      s607 <= s606;
      s608 <= s607;
      s609 <= s608;
      s610 <= s609;
      s611 <= s610;
      s612 <= s611;
      s613 <= s612;
      s614 <= s613;
      s615 <= s614;
      s616 <= s615;
      s617 <= s616;
      s618 <= s617;
      s619 <= s618;
      s620 <= s619;
      s621 <= s620;
      s622 <= s621;
      s623 <= s622;
      s624 <= s623;
      s625 <= s624;
      s626 <= s625;
      s627 <= s626;
      s628 <= s627;
      s629 <= s628;
      s630 <= s629;
      s631 <= s630;
      s632 <= s631;
      s633 <= s632;
      s634 <= s633;
      s635 <= s634;
      s636 <= s635;
      s637 <= s636;
      s638 <= s637;
      s639 <= s638;
      s640 <= s639;
      s641 <= s640;
      s642 <= s641;
      s643 <= s642;
      s644 <= s643;
      s645 <= s644;
      s646 <= s645;
      s647 <= s646;
      s648 <= s647;
      s649 <= s648;
      s650 <= s649;
      s651 <= s650;
      s652 <= s651;
      s653 <= s652;
      s654 <= s653;
      s655 <= s654;
      s656 <= s655;
      s657 <= s656;
      s658 <= s657;
      s659 <= s658;
      s660 <= s659;
      s661 <= s660;
      s662 <= s661;
      s663 <= s662;
      s664 <= s663;
      s665 <= s664;
      s666 <= s665;
      s667 <= s666;
      s668 <= s667;
      s669 <= s668;
      s670 <= s669;
      s671 <= s670;
      s672 <= s671;
      s673 <= s672;
      s674 <= s673;
      s675 <= s674;
      s676 <= s675;
      s677 <= s676;
      s678 <= s677;
      s679 <= s678;
      s680 <= s679;
      s681 <= s680;
      s682 <= s681;
      s683 <= s682;
      s684 <= s683;
      s685 <= s684;
      s686 <= s685;
      s687 <= s686;
      s688 <= s687;
      s689 <= s688;
      s690 <= s689;
      s691 <= s690;
      s692 <= s691;
      s693 <= s692;
      s694 <= s693;
      s695 <= s694;
      s696 <= s695;
      s697 <= s696;
      s698 <= s697;
      s699 <= s698;
      s700 <= s699;
      s701 <= s700;
      s702 <= s701;
      s703 <= s702;
      s704 <= s703;
      s705 <= s704;
      s706 <= s705;
      s707 <= s706;
      s708 <= s707;
      s709 <= s708;
      s710 <= s709;
      s711 <= s710;
      s712 <= s711;
      s713 <= s712;
      s714 <= s713;
      s715 <= s714;
      s716 <= s715;
      s717 <= s716;
      s718 <= s717;
      s719 <= s718;
      s720 <= s719;
      s721 <= s720;
      s722 <= s721;
      s723 <= s722;
      s724 <= s723;
      s725 <= s724;
      s726 <= s725;
      s727 <= s726;
      s728 <= s727;
      s729 <= s728;
      s730 <= s729;
      s731 <= s730;
      s732 <= s731;
      s733 <= s732;
      s734 <= s733;
      Y <= s734;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_838_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 838 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_838_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_838_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
signal s558 : std_logic_vector(33 downto 0) := (others => '0');
signal s559 : std_logic_vector(33 downto 0) := (others => '0');
signal s560 : std_logic_vector(33 downto 0) := (others => '0');
signal s561 : std_logic_vector(33 downto 0) := (others => '0');
signal s562 : std_logic_vector(33 downto 0) := (others => '0');
signal s563 : std_logic_vector(33 downto 0) := (others => '0');
signal s564 : std_logic_vector(33 downto 0) := (others => '0');
signal s565 : std_logic_vector(33 downto 0) := (others => '0');
signal s566 : std_logic_vector(33 downto 0) := (others => '0');
signal s567 : std_logic_vector(33 downto 0) := (others => '0');
signal s568 : std_logic_vector(33 downto 0) := (others => '0');
signal s569 : std_logic_vector(33 downto 0) := (others => '0');
signal s570 : std_logic_vector(33 downto 0) := (others => '0');
signal s571 : std_logic_vector(33 downto 0) := (others => '0');
signal s572 : std_logic_vector(33 downto 0) := (others => '0');
signal s573 : std_logic_vector(33 downto 0) := (others => '0');
signal s574 : std_logic_vector(33 downto 0) := (others => '0');
signal s575 : std_logic_vector(33 downto 0) := (others => '0');
signal s576 : std_logic_vector(33 downto 0) := (others => '0');
signal s577 : std_logic_vector(33 downto 0) := (others => '0');
signal s578 : std_logic_vector(33 downto 0) := (others => '0');
signal s579 : std_logic_vector(33 downto 0) := (others => '0');
signal s580 : std_logic_vector(33 downto 0) := (others => '0');
signal s581 : std_logic_vector(33 downto 0) := (others => '0');
signal s582 : std_logic_vector(33 downto 0) := (others => '0');
signal s583 : std_logic_vector(33 downto 0) := (others => '0');
signal s584 : std_logic_vector(33 downto 0) := (others => '0');
signal s585 : std_logic_vector(33 downto 0) := (others => '0');
signal s586 : std_logic_vector(33 downto 0) := (others => '0');
signal s587 : std_logic_vector(33 downto 0) := (others => '0');
signal s588 : std_logic_vector(33 downto 0) := (others => '0');
signal s589 : std_logic_vector(33 downto 0) := (others => '0');
signal s590 : std_logic_vector(33 downto 0) := (others => '0');
signal s591 : std_logic_vector(33 downto 0) := (others => '0');
signal s592 : std_logic_vector(33 downto 0) := (others => '0');
signal s593 : std_logic_vector(33 downto 0) := (others => '0');
signal s594 : std_logic_vector(33 downto 0) := (others => '0');
signal s595 : std_logic_vector(33 downto 0) := (others => '0');
signal s596 : std_logic_vector(33 downto 0) := (others => '0');
signal s597 : std_logic_vector(33 downto 0) := (others => '0');
signal s598 : std_logic_vector(33 downto 0) := (others => '0');
signal s599 : std_logic_vector(33 downto 0) := (others => '0');
signal s600 : std_logic_vector(33 downto 0) := (others => '0');
signal s601 : std_logic_vector(33 downto 0) := (others => '0');
signal s602 : std_logic_vector(33 downto 0) := (others => '0');
signal s603 : std_logic_vector(33 downto 0) := (others => '0');
signal s604 : std_logic_vector(33 downto 0) := (others => '0');
signal s605 : std_logic_vector(33 downto 0) := (others => '0');
signal s606 : std_logic_vector(33 downto 0) := (others => '0');
signal s607 : std_logic_vector(33 downto 0) := (others => '0');
signal s608 : std_logic_vector(33 downto 0) := (others => '0');
signal s609 : std_logic_vector(33 downto 0) := (others => '0');
signal s610 : std_logic_vector(33 downto 0) := (others => '0');
signal s611 : std_logic_vector(33 downto 0) := (others => '0');
signal s612 : std_logic_vector(33 downto 0) := (others => '0');
signal s613 : std_logic_vector(33 downto 0) := (others => '0');
signal s614 : std_logic_vector(33 downto 0) := (others => '0');
signal s615 : std_logic_vector(33 downto 0) := (others => '0');
signal s616 : std_logic_vector(33 downto 0) := (others => '0');
signal s617 : std_logic_vector(33 downto 0) := (others => '0');
signal s618 : std_logic_vector(33 downto 0) := (others => '0');
signal s619 : std_logic_vector(33 downto 0) := (others => '0');
signal s620 : std_logic_vector(33 downto 0) := (others => '0');
signal s621 : std_logic_vector(33 downto 0) := (others => '0');
signal s622 : std_logic_vector(33 downto 0) := (others => '0');
signal s623 : std_logic_vector(33 downto 0) := (others => '0');
signal s624 : std_logic_vector(33 downto 0) := (others => '0');
signal s625 : std_logic_vector(33 downto 0) := (others => '0');
signal s626 : std_logic_vector(33 downto 0) := (others => '0');
signal s627 : std_logic_vector(33 downto 0) := (others => '0');
signal s628 : std_logic_vector(33 downto 0) := (others => '0');
signal s629 : std_logic_vector(33 downto 0) := (others => '0');
signal s630 : std_logic_vector(33 downto 0) := (others => '0');
signal s631 : std_logic_vector(33 downto 0) := (others => '0');
signal s632 : std_logic_vector(33 downto 0) := (others => '0');
signal s633 : std_logic_vector(33 downto 0) := (others => '0');
signal s634 : std_logic_vector(33 downto 0) := (others => '0');
signal s635 : std_logic_vector(33 downto 0) := (others => '0');
signal s636 : std_logic_vector(33 downto 0) := (others => '0');
signal s637 : std_logic_vector(33 downto 0) := (others => '0');
signal s638 : std_logic_vector(33 downto 0) := (others => '0');
signal s639 : std_logic_vector(33 downto 0) := (others => '0');
signal s640 : std_logic_vector(33 downto 0) := (others => '0');
signal s641 : std_logic_vector(33 downto 0) := (others => '0');
signal s642 : std_logic_vector(33 downto 0) := (others => '0');
signal s643 : std_logic_vector(33 downto 0) := (others => '0');
signal s644 : std_logic_vector(33 downto 0) := (others => '0');
signal s645 : std_logic_vector(33 downto 0) := (others => '0');
signal s646 : std_logic_vector(33 downto 0) := (others => '0');
signal s647 : std_logic_vector(33 downto 0) := (others => '0');
signal s648 : std_logic_vector(33 downto 0) := (others => '0');
signal s649 : std_logic_vector(33 downto 0) := (others => '0');
signal s650 : std_logic_vector(33 downto 0) := (others => '0');
signal s651 : std_logic_vector(33 downto 0) := (others => '0');
signal s652 : std_logic_vector(33 downto 0) := (others => '0');
signal s653 : std_logic_vector(33 downto 0) := (others => '0');
signal s654 : std_logic_vector(33 downto 0) := (others => '0');
signal s655 : std_logic_vector(33 downto 0) := (others => '0');
signal s656 : std_logic_vector(33 downto 0) := (others => '0');
signal s657 : std_logic_vector(33 downto 0) := (others => '0');
signal s658 : std_logic_vector(33 downto 0) := (others => '0');
signal s659 : std_logic_vector(33 downto 0) := (others => '0');
signal s660 : std_logic_vector(33 downto 0) := (others => '0');
signal s661 : std_logic_vector(33 downto 0) := (others => '0');
signal s662 : std_logic_vector(33 downto 0) := (others => '0');
signal s663 : std_logic_vector(33 downto 0) := (others => '0');
signal s664 : std_logic_vector(33 downto 0) := (others => '0');
signal s665 : std_logic_vector(33 downto 0) := (others => '0');
signal s666 : std_logic_vector(33 downto 0) := (others => '0');
signal s667 : std_logic_vector(33 downto 0) := (others => '0');
signal s668 : std_logic_vector(33 downto 0) := (others => '0');
signal s669 : std_logic_vector(33 downto 0) := (others => '0');
signal s670 : std_logic_vector(33 downto 0) := (others => '0');
signal s671 : std_logic_vector(33 downto 0) := (others => '0');
signal s672 : std_logic_vector(33 downto 0) := (others => '0');
signal s673 : std_logic_vector(33 downto 0) := (others => '0');
signal s674 : std_logic_vector(33 downto 0) := (others => '0');
signal s675 : std_logic_vector(33 downto 0) := (others => '0');
signal s676 : std_logic_vector(33 downto 0) := (others => '0');
signal s677 : std_logic_vector(33 downto 0) := (others => '0');
signal s678 : std_logic_vector(33 downto 0) := (others => '0');
signal s679 : std_logic_vector(33 downto 0) := (others => '0');
signal s680 : std_logic_vector(33 downto 0) := (others => '0');
signal s681 : std_logic_vector(33 downto 0) := (others => '0');
signal s682 : std_logic_vector(33 downto 0) := (others => '0');
signal s683 : std_logic_vector(33 downto 0) := (others => '0');
signal s684 : std_logic_vector(33 downto 0) := (others => '0');
signal s685 : std_logic_vector(33 downto 0) := (others => '0');
signal s686 : std_logic_vector(33 downto 0) := (others => '0');
signal s687 : std_logic_vector(33 downto 0) := (others => '0');
signal s688 : std_logic_vector(33 downto 0) := (others => '0');
signal s689 : std_logic_vector(33 downto 0) := (others => '0');
signal s690 : std_logic_vector(33 downto 0) := (others => '0');
signal s691 : std_logic_vector(33 downto 0) := (others => '0');
signal s692 : std_logic_vector(33 downto 0) := (others => '0');
signal s693 : std_logic_vector(33 downto 0) := (others => '0');
signal s694 : std_logic_vector(33 downto 0) := (others => '0');
signal s695 : std_logic_vector(33 downto 0) := (others => '0');
signal s696 : std_logic_vector(33 downto 0) := (others => '0');
signal s697 : std_logic_vector(33 downto 0) := (others => '0');
signal s698 : std_logic_vector(33 downto 0) := (others => '0');
signal s699 : std_logic_vector(33 downto 0) := (others => '0');
signal s700 : std_logic_vector(33 downto 0) := (others => '0');
signal s701 : std_logic_vector(33 downto 0) := (others => '0');
signal s702 : std_logic_vector(33 downto 0) := (others => '0');
signal s703 : std_logic_vector(33 downto 0) := (others => '0');
signal s704 : std_logic_vector(33 downto 0) := (others => '0');
signal s705 : std_logic_vector(33 downto 0) := (others => '0');
signal s706 : std_logic_vector(33 downto 0) := (others => '0');
signal s707 : std_logic_vector(33 downto 0) := (others => '0');
signal s708 : std_logic_vector(33 downto 0) := (others => '0');
signal s709 : std_logic_vector(33 downto 0) := (others => '0');
signal s710 : std_logic_vector(33 downto 0) := (others => '0');
signal s711 : std_logic_vector(33 downto 0) := (others => '0');
signal s712 : std_logic_vector(33 downto 0) := (others => '0');
signal s713 : std_logic_vector(33 downto 0) := (others => '0');
signal s714 : std_logic_vector(33 downto 0) := (others => '0');
signal s715 : std_logic_vector(33 downto 0) := (others => '0');
signal s716 : std_logic_vector(33 downto 0) := (others => '0');
signal s717 : std_logic_vector(33 downto 0) := (others => '0');
signal s718 : std_logic_vector(33 downto 0) := (others => '0');
signal s719 : std_logic_vector(33 downto 0) := (others => '0');
signal s720 : std_logic_vector(33 downto 0) := (others => '0');
signal s721 : std_logic_vector(33 downto 0) := (others => '0');
signal s722 : std_logic_vector(33 downto 0) := (others => '0');
signal s723 : std_logic_vector(33 downto 0) := (others => '0');
signal s724 : std_logic_vector(33 downto 0) := (others => '0');
signal s725 : std_logic_vector(33 downto 0) := (others => '0');
signal s726 : std_logic_vector(33 downto 0) := (others => '0');
signal s727 : std_logic_vector(33 downto 0) := (others => '0');
signal s728 : std_logic_vector(33 downto 0) := (others => '0');
signal s729 : std_logic_vector(33 downto 0) := (others => '0');
signal s730 : std_logic_vector(33 downto 0) := (others => '0');
signal s731 : std_logic_vector(33 downto 0) := (others => '0');
signal s732 : std_logic_vector(33 downto 0) := (others => '0');
signal s733 : std_logic_vector(33 downto 0) := (others => '0');
signal s734 : std_logic_vector(33 downto 0) := (others => '0');
signal s735 : std_logic_vector(33 downto 0) := (others => '0');
signal s736 : std_logic_vector(33 downto 0) := (others => '0');
signal s737 : std_logic_vector(33 downto 0) := (others => '0');
signal s738 : std_logic_vector(33 downto 0) := (others => '0');
signal s739 : std_logic_vector(33 downto 0) := (others => '0');
signal s740 : std_logic_vector(33 downto 0) := (others => '0');
signal s741 : std_logic_vector(33 downto 0) := (others => '0');
signal s742 : std_logic_vector(33 downto 0) := (others => '0');
signal s743 : std_logic_vector(33 downto 0) := (others => '0');
signal s744 : std_logic_vector(33 downto 0) := (others => '0');
signal s745 : std_logic_vector(33 downto 0) := (others => '0');
signal s746 : std_logic_vector(33 downto 0) := (others => '0');
signal s747 : std_logic_vector(33 downto 0) := (others => '0');
signal s748 : std_logic_vector(33 downto 0) := (others => '0');
signal s749 : std_logic_vector(33 downto 0) := (others => '0');
signal s750 : std_logic_vector(33 downto 0) := (others => '0');
signal s751 : std_logic_vector(33 downto 0) := (others => '0');
signal s752 : std_logic_vector(33 downto 0) := (others => '0');
signal s753 : std_logic_vector(33 downto 0) := (others => '0');
signal s754 : std_logic_vector(33 downto 0) := (others => '0');
signal s755 : std_logic_vector(33 downto 0) := (others => '0');
signal s756 : std_logic_vector(33 downto 0) := (others => '0');
signal s757 : std_logic_vector(33 downto 0) := (others => '0');
signal s758 : std_logic_vector(33 downto 0) := (others => '0');
signal s759 : std_logic_vector(33 downto 0) := (others => '0');
signal s760 : std_logic_vector(33 downto 0) := (others => '0');
signal s761 : std_logic_vector(33 downto 0) := (others => '0');
signal s762 : std_logic_vector(33 downto 0) := (others => '0');
signal s763 : std_logic_vector(33 downto 0) := (others => '0');
signal s764 : std_logic_vector(33 downto 0) := (others => '0');
signal s765 : std_logic_vector(33 downto 0) := (others => '0');
signal s766 : std_logic_vector(33 downto 0) := (others => '0');
signal s767 : std_logic_vector(33 downto 0) := (others => '0');
signal s768 : std_logic_vector(33 downto 0) := (others => '0');
signal s769 : std_logic_vector(33 downto 0) := (others => '0');
signal s770 : std_logic_vector(33 downto 0) := (others => '0');
signal s771 : std_logic_vector(33 downto 0) := (others => '0');
signal s772 : std_logic_vector(33 downto 0) := (others => '0');
signal s773 : std_logic_vector(33 downto 0) := (others => '0');
signal s774 : std_logic_vector(33 downto 0) := (others => '0');
signal s775 : std_logic_vector(33 downto 0) := (others => '0');
signal s776 : std_logic_vector(33 downto 0) := (others => '0');
signal s777 : std_logic_vector(33 downto 0) := (others => '0');
signal s778 : std_logic_vector(33 downto 0) := (others => '0');
signal s779 : std_logic_vector(33 downto 0) := (others => '0');
signal s780 : std_logic_vector(33 downto 0) := (others => '0');
signal s781 : std_logic_vector(33 downto 0) := (others => '0');
signal s782 : std_logic_vector(33 downto 0) := (others => '0');
signal s783 : std_logic_vector(33 downto 0) := (others => '0');
signal s784 : std_logic_vector(33 downto 0) := (others => '0');
signal s785 : std_logic_vector(33 downto 0) := (others => '0');
signal s786 : std_logic_vector(33 downto 0) := (others => '0');
signal s787 : std_logic_vector(33 downto 0) := (others => '0');
signal s788 : std_logic_vector(33 downto 0) := (others => '0');
signal s789 : std_logic_vector(33 downto 0) := (others => '0');
signal s790 : std_logic_vector(33 downto 0) := (others => '0');
signal s791 : std_logic_vector(33 downto 0) := (others => '0');
signal s792 : std_logic_vector(33 downto 0) := (others => '0');
signal s793 : std_logic_vector(33 downto 0) := (others => '0');
signal s794 : std_logic_vector(33 downto 0) := (others => '0');
signal s795 : std_logic_vector(33 downto 0) := (others => '0');
signal s796 : std_logic_vector(33 downto 0) := (others => '0');
signal s797 : std_logic_vector(33 downto 0) := (others => '0');
signal s798 : std_logic_vector(33 downto 0) := (others => '0');
signal s799 : std_logic_vector(33 downto 0) := (others => '0');
signal s800 : std_logic_vector(33 downto 0) := (others => '0');
signal s801 : std_logic_vector(33 downto 0) := (others => '0');
signal s802 : std_logic_vector(33 downto 0) := (others => '0');
signal s803 : std_logic_vector(33 downto 0) := (others => '0');
signal s804 : std_logic_vector(33 downto 0) := (others => '0');
signal s805 : std_logic_vector(33 downto 0) := (others => '0');
signal s806 : std_logic_vector(33 downto 0) := (others => '0');
signal s807 : std_logic_vector(33 downto 0) := (others => '0');
signal s808 : std_logic_vector(33 downto 0) := (others => '0');
signal s809 : std_logic_vector(33 downto 0) := (others => '0');
signal s810 : std_logic_vector(33 downto 0) := (others => '0');
signal s811 : std_logic_vector(33 downto 0) := (others => '0');
signal s812 : std_logic_vector(33 downto 0) := (others => '0');
signal s813 : std_logic_vector(33 downto 0) := (others => '0');
signal s814 : std_logic_vector(33 downto 0) := (others => '0');
signal s815 : std_logic_vector(33 downto 0) := (others => '0');
signal s816 : std_logic_vector(33 downto 0) := (others => '0');
signal s817 : std_logic_vector(33 downto 0) := (others => '0');
signal s818 : std_logic_vector(33 downto 0) := (others => '0');
signal s819 : std_logic_vector(33 downto 0) := (others => '0');
signal s820 : std_logic_vector(33 downto 0) := (others => '0');
signal s821 : std_logic_vector(33 downto 0) := (others => '0');
signal s822 : std_logic_vector(33 downto 0) := (others => '0');
signal s823 : std_logic_vector(33 downto 0) := (others => '0');
signal s824 : std_logic_vector(33 downto 0) := (others => '0');
signal s825 : std_logic_vector(33 downto 0) := (others => '0');
signal s826 : std_logic_vector(33 downto 0) := (others => '0');
signal s827 : std_logic_vector(33 downto 0) := (others => '0');
signal s828 : std_logic_vector(33 downto 0) := (others => '0');
signal s829 : std_logic_vector(33 downto 0) := (others => '0');
signal s830 : std_logic_vector(33 downto 0) := (others => '0');
signal s831 : std_logic_vector(33 downto 0) := (others => '0');
signal s832 : std_logic_vector(33 downto 0) := (others => '0');
signal s833 : std_logic_vector(33 downto 0) := (others => '0');
signal s834 : std_logic_vector(33 downto 0) := (others => '0');
signal s835 : std_logic_vector(33 downto 0) := (others => '0');
signal s836 : std_logic_vector(33 downto 0) := (others => '0');
signal s837 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
      s558 <= "0000000000000000000000000000000000";
      s559 <= "0000000000000000000000000000000000";
      s560 <= "0000000000000000000000000000000000";
      s561 <= "0000000000000000000000000000000000";
      s562 <= "0000000000000000000000000000000000";
      s563 <= "0000000000000000000000000000000000";
      s564 <= "0000000000000000000000000000000000";
      s565 <= "0000000000000000000000000000000000";
      s566 <= "0000000000000000000000000000000000";
      s567 <= "0000000000000000000000000000000000";
      s568 <= "0000000000000000000000000000000000";
      s569 <= "0000000000000000000000000000000000";
      s570 <= "0000000000000000000000000000000000";
      s571 <= "0000000000000000000000000000000000";
      s572 <= "0000000000000000000000000000000000";
      s573 <= "0000000000000000000000000000000000";
      s574 <= "0000000000000000000000000000000000";
      s575 <= "0000000000000000000000000000000000";
      s576 <= "0000000000000000000000000000000000";
      s577 <= "0000000000000000000000000000000000";
      s578 <= "0000000000000000000000000000000000";
      s579 <= "0000000000000000000000000000000000";
      s580 <= "0000000000000000000000000000000000";
      s581 <= "0000000000000000000000000000000000";
      s582 <= "0000000000000000000000000000000000";
      s583 <= "0000000000000000000000000000000000";
      s584 <= "0000000000000000000000000000000000";
      s585 <= "0000000000000000000000000000000000";
      s586 <= "0000000000000000000000000000000000";
      s587 <= "0000000000000000000000000000000000";
      s588 <= "0000000000000000000000000000000000";
      s589 <= "0000000000000000000000000000000000";
      s590 <= "0000000000000000000000000000000000";
      s591 <= "0000000000000000000000000000000000";
      s592 <= "0000000000000000000000000000000000";
      s593 <= "0000000000000000000000000000000000";
      s594 <= "0000000000000000000000000000000000";
      s595 <= "0000000000000000000000000000000000";
      s596 <= "0000000000000000000000000000000000";
      s597 <= "0000000000000000000000000000000000";
      s598 <= "0000000000000000000000000000000000";
      s599 <= "0000000000000000000000000000000000";
      s600 <= "0000000000000000000000000000000000";
      s601 <= "0000000000000000000000000000000000";
      s602 <= "0000000000000000000000000000000000";
      s603 <= "0000000000000000000000000000000000";
      s604 <= "0000000000000000000000000000000000";
      s605 <= "0000000000000000000000000000000000";
      s606 <= "0000000000000000000000000000000000";
      s607 <= "0000000000000000000000000000000000";
      s608 <= "0000000000000000000000000000000000";
      s609 <= "0000000000000000000000000000000000";
      s610 <= "0000000000000000000000000000000000";
      s611 <= "0000000000000000000000000000000000";
      s612 <= "0000000000000000000000000000000000";
      s613 <= "0000000000000000000000000000000000";
      s614 <= "0000000000000000000000000000000000";
      s615 <= "0000000000000000000000000000000000";
      s616 <= "0000000000000000000000000000000000";
      s617 <= "0000000000000000000000000000000000";
      s618 <= "0000000000000000000000000000000000";
      s619 <= "0000000000000000000000000000000000";
      s620 <= "0000000000000000000000000000000000";
      s621 <= "0000000000000000000000000000000000";
      s622 <= "0000000000000000000000000000000000";
      s623 <= "0000000000000000000000000000000000";
      s624 <= "0000000000000000000000000000000000";
      s625 <= "0000000000000000000000000000000000";
      s626 <= "0000000000000000000000000000000000";
      s627 <= "0000000000000000000000000000000000";
      s628 <= "0000000000000000000000000000000000";
      s629 <= "0000000000000000000000000000000000";
      s630 <= "0000000000000000000000000000000000";
      s631 <= "0000000000000000000000000000000000";
      s632 <= "0000000000000000000000000000000000";
      s633 <= "0000000000000000000000000000000000";
      s634 <= "0000000000000000000000000000000000";
      s635 <= "0000000000000000000000000000000000";
      s636 <= "0000000000000000000000000000000000";
      s637 <= "0000000000000000000000000000000000";
      s638 <= "0000000000000000000000000000000000";
      s639 <= "0000000000000000000000000000000000";
      s640 <= "0000000000000000000000000000000000";
      s641 <= "0000000000000000000000000000000000";
      s642 <= "0000000000000000000000000000000000";
      s643 <= "0000000000000000000000000000000000";
      s644 <= "0000000000000000000000000000000000";
      s645 <= "0000000000000000000000000000000000";
      s646 <= "0000000000000000000000000000000000";
      s647 <= "0000000000000000000000000000000000";
      s648 <= "0000000000000000000000000000000000";
      s649 <= "0000000000000000000000000000000000";
      s650 <= "0000000000000000000000000000000000";
      s651 <= "0000000000000000000000000000000000";
      s652 <= "0000000000000000000000000000000000";
      s653 <= "0000000000000000000000000000000000";
      s654 <= "0000000000000000000000000000000000";
      s655 <= "0000000000000000000000000000000000";
      s656 <= "0000000000000000000000000000000000";
      s657 <= "0000000000000000000000000000000000";
      s658 <= "0000000000000000000000000000000000";
      s659 <= "0000000000000000000000000000000000";
      s660 <= "0000000000000000000000000000000000";
      s661 <= "0000000000000000000000000000000000";
      s662 <= "0000000000000000000000000000000000";
      s663 <= "0000000000000000000000000000000000";
      s664 <= "0000000000000000000000000000000000";
      s665 <= "0000000000000000000000000000000000";
      s666 <= "0000000000000000000000000000000000";
      s667 <= "0000000000000000000000000000000000";
      s668 <= "0000000000000000000000000000000000";
      s669 <= "0000000000000000000000000000000000";
      s670 <= "0000000000000000000000000000000000";
      s671 <= "0000000000000000000000000000000000";
      s672 <= "0000000000000000000000000000000000";
      s673 <= "0000000000000000000000000000000000";
      s674 <= "0000000000000000000000000000000000";
      s675 <= "0000000000000000000000000000000000";
      s676 <= "0000000000000000000000000000000000";
      s677 <= "0000000000000000000000000000000000";
      s678 <= "0000000000000000000000000000000000";
      s679 <= "0000000000000000000000000000000000";
      s680 <= "0000000000000000000000000000000000";
      s681 <= "0000000000000000000000000000000000";
      s682 <= "0000000000000000000000000000000000";
      s683 <= "0000000000000000000000000000000000";
      s684 <= "0000000000000000000000000000000000";
      s685 <= "0000000000000000000000000000000000";
      s686 <= "0000000000000000000000000000000000";
      s687 <= "0000000000000000000000000000000000";
      s688 <= "0000000000000000000000000000000000";
      s689 <= "0000000000000000000000000000000000";
      s690 <= "0000000000000000000000000000000000";
      s691 <= "0000000000000000000000000000000000";
      s692 <= "0000000000000000000000000000000000";
      s693 <= "0000000000000000000000000000000000";
      s694 <= "0000000000000000000000000000000000";
      s695 <= "0000000000000000000000000000000000";
      s696 <= "0000000000000000000000000000000000";
      s697 <= "0000000000000000000000000000000000";
      s698 <= "0000000000000000000000000000000000";
      s699 <= "0000000000000000000000000000000000";
      s700 <= "0000000000000000000000000000000000";
      s701 <= "0000000000000000000000000000000000";
      s702 <= "0000000000000000000000000000000000";
      s703 <= "0000000000000000000000000000000000";
      s704 <= "0000000000000000000000000000000000";
      s705 <= "0000000000000000000000000000000000";
      s706 <= "0000000000000000000000000000000000";
      s707 <= "0000000000000000000000000000000000";
      s708 <= "0000000000000000000000000000000000";
      s709 <= "0000000000000000000000000000000000";
      s710 <= "0000000000000000000000000000000000";
      s711 <= "0000000000000000000000000000000000";
      s712 <= "0000000000000000000000000000000000";
      s713 <= "0000000000000000000000000000000000";
      s714 <= "0000000000000000000000000000000000";
      s715 <= "0000000000000000000000000000000000";
      s716 <= "0000000000000000000000000000000000";
      s717 <= "0000000000000000000000000000000000";
      s718 <= "0000000000000000000000000000000000";
      s719 <= "0000000000000000000000000000000000";
      s720 <= "0000000000000000000000000000000000";
      s721 <= "0000000000000000000000000000000000";
      s722 <= "0000000000000000000000000000000000";
      s723 <= "0000000000000000000000000000000000";
      s724 <= "0000000000000000000000000000000000";
      s725 <= "0000000000000000000000000000000000";
      s726 <= "0000000000000000000000000000000000";
      s727 <= "0000000000000000000000000000000000";
      s728 <= "0000000000000000000000000000000000";
      s729 <= "0000000000000000000000000000000000";
      s730 <= "0000000000000000000000000000000000";
      s731 <= "0000000000000000000000000000000000";
      s732 <= "0000000000000000000000000000000000";
      s733 <= "0000000000000000000000000000000000";
      s734 <= "0000000000000000000000000000000000";
      s735 <= "0000000000000000000000000000000000";
      s736 <= "0000000000000000000000000000000000";
      s737 <= "0000000000000000000000000000000000";
      s738 <= "0000000000000000000000000000000000";
      s739 <= "0000000000000000000000000000000000";
      s740 <= "0000000000000000000000000000000000";
      s741 <= "0000000000000000000000000000000000";
      s742 <= "0000000000000000000000000000000000";
      s743 <= "0000000000000000000000000000000000";
      s744 <= "0000000000000000000000000000000000";
      s745 <= "0000000000000000000000000000000000";
      s746 <= "0000000000000000000000000000000000";
      s747 <= "0000000000000000000000000000000000";
      s748 <= "0000000000000000000000000000000000";
      s749 <= "0000000000000000000000000000000000";
      s750 <= "0000000000000000000000000000000000";
      s751 <= "0000000000000000000000000000000000";
      s752 <= "0000000000000000000000000000000000";
      s753 <= "0000000000000000000000000000000000";
      s754 <= "0000000000000000000000000000000000";
      s755 <= "0000000000000000000000000000000000";
      s756 <= "0000000000000000000000000000000000";
      s757 <= "0000000000000000000000000000000000";
      s758 <= "0000000000000000000000000000000000";
      s759 <= "0000000000000000000000000000000000";
      s760 <= "0000000000000000000000000000000000";
      s761 <= "0000000000000000000000000000000000";
      s762 <= "0000000000000000000000000000000000";
      s763 <= "0000000000000000000000000000000000";
      s764 <= "0000000000000000000000000000000000";
      s765 <= "0000000000000000000000000000000000";
      s766 <= "0000000000000000000000000000000000";
      s767 <= "0000000000000000000000000000000000";
      s768 <= "0000000000000000000000000000000000";
      s769 <= "0000000000000000000000000000000000";
      s770 <= "0000000000000000000000000000000000";
      s771 <= "0000000000000000000000000000000000";
      s772 <= "0000000000000000000000000000000000";
      s773 <= "0000000000000000000000000000000000";
      s774 <= "0000000000000000000000000000000000";
      s775 <= "0000000000000000000000000000000000";
      s776 <= "0000000000000000000000000000000000";
      s777 <= "0000000000000000000000000000000000";
      s778 <= "0000000000000000000000000000000000";
      s779 <= "0000000000000000000000000000000000";
      s780 <= "0000000000000000000000000000000000";
      s781 <= "0000000000000000000000000000000000";
      s782 <= "0000000000000000000000000000000000";
      s783 <= "0000000000000000000000000000000000";
      s784 <= "0000000000000000000000000000000000";
      s785 <= "0000000000000000000000000000000000";
      s786 <= "0000000000000000000000000000000000";
      s787 <= "0000000000000000000000000000000000";
      s788 <= "0000000000000000000000000000000000";
      s789 <= "0000000000000000000000000000000000";
      s790 <= "0000000000000000000000000000000000";
      s791 <= "0000000000000000000000000000000000";
      s792 <= "0000000000000000000000000000000000";
      s793 <= "0000000000000000000000000000000000";
      s794 <= "0000000000000000000000000000000000";
      s795 <= "0000000000000000000000000000000000";
      s796 <= "0000000000000000000000000000000000";
      s797 <= "0000000000000000000000000000000000";
      s798 <= "0000000000000000000000000000000000";
      s799 <= "0000000000000000000000000000000000";
      s800 <= "0000000000000000000000000000000000";
      s801 <= "0000000000000000000000000000000000";
      s802 <= "0000000000000000000000000000000000";
      s803 <= "0000000000000000000000000000000000";
      s804 <= "0000000000000000000000000000000000";
      s805 <= "0000000000000000000000000000000000";
      s806 <= "0000000000000000000000000000000000";
      s807 <= "0000000000000000000000000000000000";
      s808 <= "0000000000000000000000000000000000";
      s809 <= "0000000000000000000000000000000000";
      s810 <= "0000000000000000000000000000000000";
      s811 <= "0000000000000000000000000000000000";
      s812 <= "0000000000000000000000000000000000";
      s813 <= "0000000000000000000000000000000000";
      s814 <= "0000000000000000000000000000000000";
      s815 <= "0000000000000000000000000000000000";
      s816 <= "0000000000000000000000000000000000";
      s817 <= "0000000000000000000000000000000000";
      s818 <= "0000000000000000000000000000000000";
      s819 <= "0000000000000000000000000000000000";
      s820 <= "0000000000000000000000000000000000";
      s821 <= "0000000000000000000000000000000000";
      s822 <= "0000000000000000000000000000000000";
      s823 <= "0000000000000000000000000000000000";
      s824 <= "0000000000000000000000000000000000";
      s825 <= "0000000000000000000000000000000000";
      s826 <= "0000000000000000000000000000000000";
      s827 <= "0000000000000000000000000000000000";
      s828 <= "0000000000000000000000000000000000";
      s829 <= "0000000000000000000000000000000000";
      s830 <= "0000000000000000000000000000000000";
      s831 <= "0000000000000000000000000000000000";
      s832 <= "0000000000000000000000000000000000";
      s833 <= "0000000000000000000000000000000000";
      s834 <= "0000000000000000000000000000000000";
      s835 <= "0000000000000000000000000000000000";
      s836 <= "0000000000000000000000000000000000";
      s837 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      s558 <= s557;
      s559 <= s558;
      s560 <= s559;
      s561 <= s560;
      s562 <= s561;
      s563 <= s562;
      s564 <= s563;
      s565 <= s564;
      s566 <= s565;
      s567 <= s566;
      s568 <= s567;
      s569 <= s568;
      s570 <= s569;
      s571 <= s570;
      s572 <= s571;
      s573 <= s572;
      s574 <= s573;
      s575 <= s574;
      s576 <= s575;
      s577 <= s576;
      s578 <= s577;
      s579 <= s578;
      s580 <= s579;
      s581 <= s580;
      s582 <= s581;
      s583 <= s582;
      s584 <= s583;
      s585 <= s584;
      s586 <= s585;
      s587 <= s586;
      s588 <= s587;
      s589 <= s588;
      s590 <= s589;
      s591 <= s590;
      s592 <= s591;
      s593 <= s592;
      s594 <= s593;
      s595 <= s594;
      s596 <= s595;
      s597 <= s596;
      s598 <= s597;
      s599 <= s598;
      s600 <= s599;
      s601 <= s600;
      s602 <= s601;
      s603 <= s602;
      s604 <= s603;
      s605 <= s604;
      s606 <= s605;
      s607 <= s606;
      s608 <= s607;
      s609 <= s608;
      s610 <= s609;
      s611 <= s610;
      s612 <= s611;
      s613 <= s612;
      s614 <= s613;
      s615 <= s614;
      s616 <= s615;
      s617 <= s616;
      s618 <= s617;
      s619 <= s618;
      s620 <= s619;
      s621 <= s620;
      s622 <= s621;
      s623 <= s622;
      s624 <= s623;
      s625 <= s624;
      s626 <= s625;
      s627 <= s626;
      s628 <= s627;
      s629 <= s628;
      s630 <= s629;
      s631 <= s630;
      s632 <= s631;
      s633 <= s632;
      s634 <= s633;
      s635 <= s634;
      s636 <= s635;
      s637 <= s636;
      s638 <= s637;
      s639 <= s638;
      s640 <= s639;
      s641 <= s640;
      s642 <= s641;
      s643 <= s642;
      s644 <= s643;
      s645 <= s644;
      s646 <= s645;
      s647 <= s646;
      s648 <= s647;
      s649 <= s648;
      s650 <= s649;
      s651 <= s650;
      s652 <= s651;
      s653 <= s652;
      s654 <= s653;
      s655 <= s654;
      s656 <= s655;
      s657 <= s656;
      s658 <= s657;
      s659 <= s658;
      s660 <= s659;
      s661 <= s660;
      s662 <= s661;
      s663 <= s662;
      s664 <= s663;
      s665 <= s664;
      s666 <= s665;
      s667 <= s666;
      s668 <= s667;
      s669 <= s668;
      s670 <= s669;
      s671 <= s670;
      s672 <= s671;
      s673 <= s672;
      s674 <= s673;
      s675 <= s674;
      s676 <= s675;
      s677 <= s676;
      s678 <= s677;
      s679 <= s678;
      s680 <= s679;
      s681 <= s680;
      s682 <= s681;
      s683 <= s682;
      s684 <= s683;
      s685 <= s684;
      s686 <= s685;
      s687 <= s686;
      s688 <= s687;
      s689 <= s688;
      s690 <= s689;
      s691 <= s690;
      s692 <= s691;
      s693 <= s692;
      s694 <= s693;
      s695 <= s694;
      s696 <= s695;
      s697 <= s696;
      s698 <= s697;
      s699 <= s698;
      s700 <= s699;
      s701 <= s700;
      s702 <= s701;
      s703 <= s702;
      s704 <= s703;
      s705 <= s704;
      s706 <= s705;
      s707 <= s706;
      s708 <= s707;
      s709 <= s708;
      s710 <= s709;
      s711 <= s710;
      s712 <= s711;
      s713 <= s712;
      s714 <= s713;
      s715 <= s714;
      s716 <= s715;
      s717 <= s716;
      s718 <= s717;
      s719 <= s718;
      s720 <= s719;
      s721 <= s720;
      s722 <= s721;
      s723 <= s722;
      s724 <= s723;
      s725 <= s724;
      s726 <= s725;
      s727 <= s726;
      s728 <= s727;
      s729 <= s728;
      s730 <= s729;
      s731 <= s730;
      s732 <= s731;
      s733 <= s732;
      s734 <= s733;
      s735 <= s734;
      s736 <= s735;
      s737 <= s736;
      s738 <= s737;
      s739 <= s738;
      s740 <= s739;
      s741 <= s740;
      s742 <= s741;
      s743 <= s742;
      s744 <= s743;
      s745 <= s744;
      s746 <= s745;
      s747 <= s746;
      s748 <= s747;
      s749 <= s748;
      s750 <= s749;
      s751 <= s750;
      s752 <= s751;
      s753 <= s752;
      s754 <= s753;
      s755 <= s754;
      s756 <= s755;
      s757 <= s756;
      s758 <= s757;
      s759 <= s758;
      s760 <= s759;
      s761 <= s760;
      s762 <= s761;
      s763 <= s762;
      s764 <= s763;
      s765 <= s764;
      s766 <= s765;
      s767 <= s766;
      s768 <= s767;
      s769 <= s768;
      s770 <= s769;
      s771 <= s770;
      s772 <= s771;
      s773 <= s772;
      s774 <= s773;
      s775 <= s774;
      s776 <= s775;
      s777 <= s776;
      s778 <= s777;
      s779 <= s778;
      s780 <= s779;
      s781 <= s780;
      s782 <= s781;
      s783 <= s782;
      s784 <= s783;
      s785 <= s784;
      s786 <= s785;
      s787 <= s786;
      s788 <= s787;
      s789 <= s788;
      s790 <= s789;
      s791 <= s790;
      s792 <= s791;
      s793 <= s792;
      s794 <= s793;
      s795 <= s794;
      s796 <= s795;
      s797 <= s796;
      s798 <= s797;
      s799 <= s798;
      s800 <= s799;
      s801 <= s800;
      s802 <= s801;
      s803 <= s802;
      s804 <= s803;
      s805 <= s804;
      s806 <= s805;
      s807 <= s806;
      s808 <= s807;
      s809 <= s808;
      s810 <= s809;
      s811 <= s810;
      s812 <= s811;
      s813 <= s812;
      s814 <= s813;
      s815 <= s814;
      s816 <= s815;
      s817 <= s816;
      s818 <= s817;
      s819 <= s818;
      s820 <= s819;
      s821 <= s820;
      s822 <= s821;
      s823 <= s822;
      s824 <= s823;
      s825 <= s824;
      s826 <= s825;
      s827 <= s826;
      s828 <= s827;
      s829 <= s828;
      s830 <= s829;
      s831 <= s830;
      s832 <= s831;
      s833 <= s832;
      s834 <= s833;
      s835 <= s834;
      s836 <= s835;
      s837 <= s836;
      Y <= s837;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_946_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 946 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_946_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_946_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
signal s558 : std_logic_vector(33 downto 0) := (others => '0');
signal s559 : std_logic_vector(33 downto 0) := (others => '0');
signal s560 : std_logic_vector(33 downto 0) := (others => '0');
signal s561 : std_logic_vector(33 downto 0) := (others => '0');
signal s562 : std_logic_vector(33 downto 0) := (others => '0');
signal s563 : std_logic_vector(33 downto 0) := (others => '0');
signal s564 : std_logic_vector(33 downto 0) := (others => '0');
signal s565 : std_logic_vector(33 downto 0) := (others => '0');
signal s566 : std_logic_vector(33 downto 0) := (others => '0');
signal s567 : std_logic_vector(33 downto 0) := (others => '0');
signal s568 : std_logic_vector(33 downto 0) := (others => '0');
signal s569 : std_logic_vector(33 downto 0) := (others => '0');
signal s570 : std_logic_vector(33 downto 0) := (others => '0');
signal s571 : std_logic_vector(33 downto 0) := (others => '0');
signal s572 : std_logic_vector(33 downto 0) := (others => '0');
signal s573 : std_logic_vector(33 downto 0) := (others => '0');
signal s574 : std_logic_vector(33 downto 0) := (others => '0');
signal s575 : std_logic_vector(33 downto 0) := (others => '0');
signal s576 : std_logic_vector(33 downto 0) := (others => '0');
signal s577 : std_logic_vector(33 downto 0) := (others => '0');
signal s578 : std_logic_vector(33 downto 0) := (others => '0');
signal s579 : std_logic_vector(33 downto 0) := (others => '0');
signal s580 : std_logic_vector(33 downto 0) := (others => '0');
signal s581 : std_logic_vector(33 downto 0) := (others => '0');
signal s582 : std_logic_vector(33 downto 0) := (others => '0');
signal s583 : std_logic_vector(33 downto 0) := (others => '0');
signal s584 : std_logic_vector(33 downto 0) := (others => '0');
signal s585 : std_logic_vector(33 downto 0) := (others => '0');
signal s586 : std_logic_vector(33 downto 0) := (others => '0');
signal s587 : std_logic_vector(33 downto 0) := (others => '0');
signal s588 : std_logic_vector(33 downto 0) := (others => '0');
signal s589 : std_logic_vector(33 downto 0) := (others => '0');
signal s590 : std_logic_vector(33 downto 0) := (others => '0');
signal s591 : std_logic_vector(33 downto 0) := (others => '0');
signal s592 : std_logic_vector(33 downto 0) := (others => '0');
signal s593 : std_logic_vector(33 downto 0) := (others => '0');
signal s594 : std_logic_vector(33 downto 0) := (others => '0');
signal s595 : std_logic_vector(33 downto 0) := (others => '0');
signal s596 : std_logic_vector(33 downto 0) := (others => '0');
signal s597 : std_logic_vector(33 downto 0) := (others => '0');
signal s598 : std_logic_vector(33 downto 0) := (others => '0');
signal s599 : std_logic_vector(33 downto 0) := (others => '0');
signal s600 : std_logic_vector(33 downto 0) := (others => '0');
signal s601 : std_logic_vector(33 downto 0) := (others => '0');
signal s602 : std_logic_vector(33 downto 0) := (others => '0');
signal s603 : std_logic_vector(33 downto 0) := (others => '0');
signal s604 : std_logic_vector(33 downto 0) := (others => '0');
signal s605 : std_logic_vector(33 downto 0) := (others => '0');
signal s606 : std_logic_vector(33 downto 0) := (others => '0');
signal s607 : std_logic_vector(33 downto 0) := (others => '0');
signal s608 : std_logic_vector(33 downto 0) := (others => '0');
signal s609 : std_logic_vector(33 downto 0) := (others => '0');
signal s610 : std_logic_vector(33 downto 0) := (others => '0');
signal s611 : std_logic_vector(33 downto 0) := (others => '0');
signal s612 : std_logic_vector(33 downto 0) := (others => '0');
signal s613 : std_logic_vector(33 downto 0) := (others => '0');
signal s614 : std_logic_vector(33 downto 0) := (others => '0');
signal s615 : std_logic_vector(33 downto 0) := (others => '0');
signal s616 : std_logic_vector(33 downto 0) := (others => '0');
signal s617 : std_logic_vector(33 downto 0) := (others => '0');
signal s618 : std_logic_vector(33 downto 0) := (others => '0');
signal s619 : std_logic_vector(33 downto 0) := (others => '0');
signal s620 : std_logic_vector(33 downto 0) := (others => '0');
signal s621 : std_logic_vector(33 downto 0) := (others => '0');
signal s622 : std_logic_vector(33 downto 0) := (others => '0');
signal s623 : std_logic_vector(33 downto 0) := (others => '0');
signal s624 : std_logic_vector(33 downto 0) := (others => '0');
signal s625 : std_logic_vector(33 downto 0) := (others => '0');
signal s626 : std_logic_vector(33 downto 0) := (others => '0');
signal s627 : std_logic_vector(33 downto 0) := (others => '0');
signal s628 : std_logic_vector(33 downto 0) := (others => '0');
signal s629 : std_logic_vector(33 downto 0) := (others => '0');
signal s630 : std_logic_vector(33 downto 0) := (others => '0');
signal s631 : std_logic_vector(33 downto 0) := (others => '0');
signal s632 : std_logic_vector(33 downto 0) := (others => '0');
signal s633 : std_logic_vector(33 downto 0) := (others => '0');
signal s634 : std_logic_vector(33 downto 0) := (others => '0');
signal s635 : std_logic_vector(33 downto 0) := (others => '0');
signal s636 : std_logic_vector(33 downto 0) := (others => '0');
signal s637 : std_logic_vector(33 downto 0) := (others => '0');
signal s638 : std_logic_vector(33 downto 0) := (others => '0');
signal s639 : std_logic_vector(33 downto 0) := (others => '0');
signal s640 : std_logic_vector(33 downto 0) := (others => '0');
signal s641 : std_logic_vector(33 downto 0) := (others => '0');
signal s642 : std_logic_vector(33 downto 0) := (others => '0');
signal s643 : std_logic_vector(33 downto 0) := (others => '0');
signal s644 : std_logic_vector(33 downto 0) := (others => '0');
signal s645 : std_logic_vector(33 downto 0) := (others => '0');
signal s646 : std_logic_vector(33 downto 0) := (others => '0');
signal s647 : std_logic_vector(33 downto 0) := (others => '0');
signal s648 : std_logic_vector(33 downto 0) := (others => '0');
signal s649 : std_logic_vector(33 downto 0) := (others => '0');
signal s650 : std_logic_vector(33 downto 0) := (others => '0');
signal s651 : std_logic_vector(33 downto 0) := (others => '0');
signal s652 : std_logic_vector(33 downto 0) := (others => '0');
signal s653 : std_logic_vector(33 downto 0) := (others => '0');
signal s654 : std_logic_vector(33 downto 0) := (others => '0');
signal s655 : std_logic_vector(33 downto 0) := (others => '0');
signal s656 : std_logic_vector(33 downto 0) := (others => '0');
signal s657 : std_logic_vector(33 downto 0) := (others => '0');
signal s658 : std_logic_vector(33 downto 0) := (others => '0');
signal s659 : std_logic_vector(33 downto 0) := (others => '0');
signal s660 : std_logic_vector(33 downto 0) := (others => '0');
signal s661 : std_logic_vector(33 downto 0) := (others => '0');
signal s662 : std_logic_vector(33 downto 0) := (others => '0');
signal s663 : std_logic_vector(33 downto 0) := (others => '0');
signal s664 : std_logic_vector(33 downto 0) := (others => '0');
signal s665 : std_logic_vector(33 downto 0) := (others => '0');
signal s666 : std_logic_vector(33 downto 0) := (others => '0');
signal s667 : std_logic_vector(33 downto 0) := (others => '0');
signal s668 : std_logic_vector(33 downto 0) := (others => '0');
signal s669 : std_logic_vector(33 downto 0) := (others => '0');
signal s670 : std_logic_vector(33 downto 0) := (others => '0');
signal s671 : std_logic_vector(33 downto 0) := (others => '0');
signal s672 : std_logic_vector(33 downto 0) := (others => '0');
signal s673 : std_logic_vector(33 downto 0) := (others => '0');
signal s674 : std_logic_vector(33 downto 0) := (others => '0');
signal s675 : std_logic_vector(33 downto 0) := (others => '0');
signal s676 : std_logic_vector(33 downto 0) := (others => '0');
signal s677 : std_logic_vector(33 downto 0) := (others => '0');
signal s678 : std_logic_vector(33 downto 0) := (others => '0');
signal s679 : std_logic_vector(33 downto 0) := (others => '0');
signal s680 : std_logic_vector(33 downto 0) := (others => '0');
signal s681 : std_logic_vector(33 downto 0) := (others => '0');
signal s682 : std_logic_vector(33 downto 0) := (others => '0');
signal s683 : std_logic_vector(33 downto 0) := (others => '0');
signal s684 : std_logic_vector(33 downto 0) := (others => '0');
signal s685 : std_logic_vector(33 downto 0) := (others => '0');
signal s686 : std_logic_vector(33 downto 0) := (others => '0');
signal s687 : std_logic_vector(33 downto 0) := (others => '0');
signal s688 : std_logic_vector(33 downto 0) := (others => '0');
signal s689 : std_logic_vector(33 downto 0) := (others => '0');
signal s690 : std_logic_vector(33 downto 0) := (others => '0');
signal s691 : std_logic_vector(33 downto 0) := (others => '0');
signal s692 : std_logic_vector(33 downto 0) := (others => '0');
signal s693 : std_logic_vector(33 downto 0) := (others => '0');
signal s694 : std_logic_vector(33 downto 0) := (others => '0');
signal s695 : std_logic_vector(33 downto 0) := (others => '0');
signal s696 : std_logic_vector(33 downto 0) := (others => '0');
signal s697 : std_logic_vector(33 downto 0) := (others => '0');
signal s698 : std_logic_vector(33 downto 0) := (others => '0');
signal s699 : std_logic_vector(33 downto 0) := (others => '0');
signal s700 : std_logic_vector(33 downto 0) := (others => '0');
signal s701 : std_logic_vector(33 downto 0) := (others => '0');
signal s702 : std_logic_vector(33 downto 0) := (others => '0');
signal s703 : std_logic_vector(33 downto 0) := (others => '0');
signal s704 : std_logic_vector(33 downto 0) := (others => '0');
signal s705 : std_logic_vector(33 downto 0) := (others => '0');
signal s706 : std_logic_vector(33 downto 0) := (others => '0');
signal s707 : std_logic_vector(33 downto 0) := (others => '0');
signal s708 : std_logic_vector(33 downto 0) := (others => '0');
signal s709 : std_logic_vector(33 downto 0) := (others => '0');
signal s710 : std_logic_vector(33 downto 0) := (others => '0');
signal s711 : std_logic_vector(33 downto 0) := (others => '0');
signal s712 : std_logic_vector(33 downto 0) := (others => '0');
signal s713 : std_logic_vector(33 downto 0) := (others => '0');
signal s714 : std_logic_vector(33 downto 0) := (others => '0');
signal s715 : std_logic_vector(33 downto 0) := (others => '0');
signal s716 : std_logic_vector(33 downto 0) := (others => '0');
signal s717 : std_logic_vector(33 downto 0) := (others => '0');
signal s718 : std_logic_vector(33 downto 0) := (others => '0');
signal s719 : std_logic_vector(33 downto 0) := (others => '0');
signal s720 : std_logic_vector(33 downto 0) := (others => '0');
signal s721 : std_logic_vector(33 downto 0) := (others => '0');
signal s722 : std_logic_vector(33 downto 0) := (others => '0');
signal s723 : std_logic_vector(33 downto 0) := (others => '0');
signal s724 : std_logic_vector(33 downto 0) := (others => '0');
signal s725 : std_logic_vector(33 downto 0) := (others => '0');
signal s726 : std_logic_vector(33 downto 0) := (others => '0');
signal s727 : std_logic_vector(33 downto 0) := (others => '0');
signal s728 : std_logic_vector(33 downto 0) := (others => '0');
signal s729 : std_logic_vector(33 downto 0) := (others => '0');
signal s730 : std_logic_vector(33 downto 0) := (others => '0');
signal s731 : std_logic_vector(33 downto 0) := (others => '0');
signal s732 : std_logic_vector(33 downto 0) := (others => '0');
signal s733 : std_logic_vector(33 downto 0) := (others => '0');
signal s734 : std_logic_vector(33 downto 0) := (others => '0');
signal s735 : std_logic_vector(33 downto 0) := (others => '0');
signal s736 : std_logic_vector(33 downto 0) := (others => '0');
signal s737 : std_logic_vector(33 downto 0) := (others => '0');
signal s738 : std_logic_vector(33 downto 0) := (others => '0');
signal s739 : std_logic_vector(33 downto 0) := (others => '0');
signal s740 : std_logic_vector(33 downto 0) := (others => '0');
signal s741 : std_logic_vector(33 downto 0) := (others => '0');
signal s742 : std_logic_vector(33 downto 0) := (others => '0');
signal s743 : std_logic_vector(33 downto 0) := (others => '0');
signal s744 : std_logic_vector(33 downto 0) := (others => '0');
signal s745 : std_logic_vector(33 downto 0) := (others => '0');
signal s746 : std_logic_vector(33 downto 0) := (others => '0');
signal s747 : std_logic_vector(33 downto 0) := (others => '0');
signal s748 : std_logic_vector(33 downto 0) := (others => '0');
signal s749 : std_logic_vector(33 downto 0) := (others => '0');
signal s750 : std_logic_vector(33 downto 0) := (others => '0');
signal s751 : std_logic_vector(33 downto 0) := (others => '0');
signal s752 : std_logic_vector(33 downto 0) := (others => '0');
signal s753 : std_logic_vector(33 downto 0) := (others => '0');
signal s754 : std_logic_vector(33 downto 0) := (others => '0');
signal s755 : std_logic_vector(33 downto 0) := (others => '0');
signal s756 : std_logic_vector(33 downto 0) := (others => '0');
signal s757 : std_logic_vector(33 downto 0) := (others => '0');
signal s758 : std_logic_vector(33 downto 0) := (others => '0');
signal s759 : std_logic_vector(33 downto 0) := (others => '0');
signal s760 : std_logic_vector(33 downto 0) := (others => '0');
signal s761 : std_logic_vector(33 downto 0) := (others => '0');
signal s762 : std_logic_vector(33 downto 0) := (others => '0');
signal s763 : std_logic_vector(33 downto 0) := (others => '0');
signal s764 : std_logic_vector(33 downto 0) := (others => '0');
signal s765 : std_logic_vector(33 downto 0) := (others => '0');
signal s766 : std_logic_vector(33 downto 0) := (others => '0');
signal s767 : std_logic_vector(33 downto 0) := (others => '0');
signal s768 : std_logic_vector(33 downto 0) := (others => '0');
signal s769 : std_logic_vector(33 downto 0) := (others => '0');
signal s770 : std_logic_vector(33 downto 0) := (others => '0');
signal s771 : std_logic_vector(33 downto 0) := (others => '0');
signal s772 : std_logic_vector(33 downto 0) := (others => '0');
signal s773 : std_logic_vector(33 downto 0) := (others => '0');
signal s774 : std_logic_vector(33 downto 0) := (others => '0');
signal s775 : std_logic_vector(33 downto 0) := (others => '0');
signal s776 : std_logic_vector(33 downto 0) := (others => '0');
signal s777 : std_logic_vector(33 downto 0) := (others => '0');
signal s778 : std_logic_vector(33 downto 0) := (others => '0');
signal s779 : std_logic_vector(33 downto 0) := (others => '0');
signal s780 : std_logic_vector(33 downto 0) := (others => '0');
signal s781 : std_logic_vector(33 downto 0) := (others => '0');
signal s782 : std_logic_vector(33 downto 0) := (others => '0');
signal s783 : std_logic_vector(33 downto 0) := (others => '0');
signal s784 : std_logic_vector(33 downto 0) := (others => '0');
signal s785 : std_logic_vector(33 downto 0) := (others => '0');
signal s786 : std_logic_vector(33 downto 0) := (others => '0');
signal s787 : std_logic_vector(33 downto 0) := (others => '0');
signal s788 : std_logic_vector(33 downto 0) := (others => '0');
signal s789 : std_logic_vector(33 downto 0) := (others => '0');
signal s790 : std_logic_vector(33 downto 0) := (others => '0');
signal s791 : std_logic_vector(33 downto 0) := (others => '0');
signal s792 : std_logic_vector(33 downto 0) := (others => '0');
signal s793 : std_logic_vector(33 downto 0) := (others => '0');
signal s794 : std_logic_vector(33 downto 0) := (others => '0');
signal s795 : std_logic_vector(33 downto 0) := (others => '0');
signal s796 : std_logic_vector(33 downto 0) := (others => '0');
signal s797 : std_logic_vector(33 downto 0) := (others => '0');
signal s798 : std_logic_vector(33 downto 0) := (others => '0');
signal s799 : std_logic_vector(33 downto 0) := (others => '0');
signal s800 : std_logic_vector(33 downto 0) := (others => '0');
signal s801 : std_logic_vector(33 downto 0) := (others => '0');
signal s802 : std_logic_vector(33 downto 0) := (others => '0');
signal s803 : std_logic_vector(33 downto 0) := (others => '0');
signal s804 : std_logic_vector(33 downto 0) := (others => '0');
signal s805 : std_logic_vector(33 downto 0) := (others => '0');
signal s806 : std_logic_vector(33 downto 0) := (others => '0');
signal s807 : std_logic_vector(33 downto 0) := (others => '0');
signal s808 : std_logic_vector(33 downto 0) := (others => '0');
signal s809 : std_logic_vector(33 downto 0) := (others => '0');
signal s810 : std_logic_vector(33 downto 0) := (others => '0');
signal s811 : std_logic_vector(33 downto 0) := (others => '0');
signal s812 : std_logic_vector(33 downto 0) := (others => '0');
signal s813 : std_logic_vector(33 downto 0) := (others => '0');
signal s814 : std_logic_vector(33 downto 0) := (others => '0');
signal s815 : std_logic_vector(33 downto 0) := (others => '0');
signal s816 : std_logic_vector(33 downto 0) := (others => '0');
signal s817 : std_logic_vector(33 downto 0) := (others => '0');
signal s818 : std_logic_vector(33 downto 0) := (others => '0');
signal s819 : std_logic_vector(33 downto 0) := (others => '0');
signal s820 : std_logic_vector(33 downto 0) := (others => '0');
signal s821 : std_logic_vector(33 downto 0) := (others => '0');
signal s822 : std_logic_vector(33 downto 0) := (others => '0');
signal s823 : std_logic_vector(33 downto 0) := (others => '0');
signal s824 : std_logic_vector(33 downto 0) := (others => '0');
signal s825 : std_logic_vector(33 downto 0) := (others => '0');
signal s826 : std_logic_vector(33 downto 0) := (others => '0');
signal s827 : std_logic_vector(33 downto 0) := (others => '0');
signal s828 : std_logic_vector(33 downto 0) := (others => '0');
signal s829 : std_logic_vector(33 downto 0) := (others => '0');
signal s830 : std_logic_vector(33 downto 0) := (others => '0');
signal s831 : std_logic_vector(33 downto 0) := (others => '0');
signal s832 : std_logic_vector(33 downto 0) := (others => '0');
signal s833 : std_logic_vector(33 downto 0) := (others => '0');
signal s834 : std_logic_vector(33 downto 0) := (others => '0');
signal s835 : std_logic_vector(33 downto 0) := (others => '0');
signal s836 : std_logic_vector(33 downto 0) := (others => '0');
signal s837 : std_logic_vector(33 downto 0) := (others => '0');
signal s838 : std_logic_vector(33 downto 0) := (others => '0');
signal s839 : std_logic_vector(33 downto 0) := (others => '0');
signal s840 : std_logic_vector(33 downto 0) := (others => '0');
signal s841 : std_logic_vector(33 downto 0) := (others => '0');
signal s842 : std_logic_vector(33 downto 0) := (others => '0');
signal s843 : std_logic_vector(33 downto 0) := (others => '0');
signal s844 : std_logic_vector(33 downto 0) := (others => '0');
signal s845 : std_logic_vector(33 downto 0) := (others => '0');
signal s846 : std_logic_vector(33 downto 0) := (others => '0');
signal s847 : std_logic_vector(33 downto 0) := (others => '0');
signal s848 : std_logic_vector(33 downto 0) := (others => '0');
signal s849 : std_logic_vector(33 downto 0) := (others => '0');
signal s850 : std_logic_vector(33 downto 0) := (others => '0');
signal s851 : std_logic_vector(33 downto 0) := (others => '0');
signal s852 : std_logic_vector(33 downto 0) := (others => '0');
signal s853 : std_logic_vector(33 downto 0) := (others => '0');
signal s854 : std_logic_vector(33 downto 0) := (others => '0');
signal s855 : std_logic_vector(33 downto 0) := (others => '0');
signal s856 : std_logic_vector(33 downto 0) := (others => '0');
signal s857 : std_logic_vector(33 downto 0) := (others => '0');
signal s858 : std_logic_vector(33 downto 0) := (others => '0');
signal s859 : std_logic_vector(33 downto 0) := (others => '0');
signal s860 : std_logic_vector(33 downto 0) := (others => '0');
signal s861 : std_logic_vector(33 downto 0) := (others => '0');
signal s862 : std_logic_vector(33 downto 0) := (others => '0');
signal s863 : std_logic_vector(33 downto 0) := (others => '0');
signal s864 : std_logic_vector(33 downto 0) := (others => '0');
signal s865 : std_logic_vector(33 downto 0) := (others => '0');
signal s866 : std_logic_vector(33 downto 0) := (others => '0');
signal s867 : std_logic_vector(33 downto 0) := (others => '0');
signal s868 : std_logic_vector(33 downto 0) := (others => '0');
signal s869 : std_logic_vector(33 downto 0) := (others => '0');
signal s870 : std_logic_vector(33 downto 0) := (others => '0');
signal s871 : std_logic_vector(33 downto 0) := (others => '0');
signal s872 : std_logic_vector(33 downto 0) := (others => '0');
signal s873 : std_logic_vector(33 downto 0) := (others => '0');
signal s874 : std_logic_vector(33 downto 0) := (others => '0');
signal s875 : std_logic_vector(33 downto 0) := (others => '0');
signal s876 : std_logic_vector(33 downto 0) := (others => '0');
signal s877 : std_logic_vector(33 downto 0) := (others => '0');
signal s878 : std_logic_vector(33 downto 0) := (others => '0');
signal s879 : std_logic_vector(33 downto 0) := (others => '0');
signal s880 : std_logic_vector(33 downto 0) := (others => '0');
signal s881 : std_logic_vector(33 downto 0) := (others => '0');
signal s882 : std_logic_vector(33 downto 0) := (others => '0');
signal s883 : std_logic_vector(33 downto 0) := (others => '0');
signal s884 : std_logic_vector(33 downto 0) := (others => '0');
signal s885 : std_logic_vector(33 downto 0) := (others => '0');
signal s886 : std_logic_vector(33 downto 0) := (others => '0');
signal s887 : std_logic_vector(33 downto 0) := (others => '0');
signal s888 : std_logic_vector(33 downto 0) := (others => '0');
signal s889 : std_logic_vector(33 downto 0) := (others => '0');
signal s890 : std_logic_vector(33 downto 0) := (others => '0');
signal s891 : std_logic_vector(33 downto 0) := (others => '0');
signal s892 : std_logic_vector(33 downto 0) := (others => '0');
signal s893 : std_logic_vector(33 downto 0) := (others => '0');
signal s894 : std_logic_vector(33 downto 0) := (others => '0');
signal s895 : std_logic_vector(33 downto 0) := (others => '0');
signal s896 : std_logic_vector(33 downto 0) := (others => '0');
signal s897 : std_logic_vector(33 downto 0) := (others => '0');
signal s898 : std_logic_vector(33 downto 0) := (others => '0');
signal s899 : std_logic_vector(33 downto 0) := (others => '0');
signal s900 : std_logic_vector(33 downto 0) := (others => '0');
signal s901 : std_logic_vector(33 downto 0) := (others => '0');
signal s902 : std_logic_vector(33 downto 0) := (others => '0');
signal s903 : std_logic_vector(33 downto 0) := (others => '0');
signal s904 : std_logic_vector(33 downto 0) := (others => '0');
signal s905 : std_logic_vector(33 downto 0) := (others => '0');
signal s906 : std_logic_vector(33 downto 0) := (others => '0');
signal s907 : std_logic_vector(33 downto 0) := (others => '0');
signal s908 : std_logic_vector(33 downto 0) := (others => '0');
signal s909 : std_logic_vector(33 downto 0) := (others => '0');
signal s910 : std_logic_vector(33 downto 0) := (others => '0');
signal s911 : std_logic_vector(33 downto 0) := (others => '0');
signal s912 : std_logic_vector(33 downto 0) := (others => '0');
signal s913 : std_logic_vector(33 downto 0) := (others => '0');
signal s914 : std_logic_vector(33 downto 0) := (others => '0');
signal s915 : std_logic_vector(33 downto 0) := (others => '0');
signal s916 : std_logic_vector(33 downto 0) := (others => '0');
signal s917 : std_logic_vector(33 downto 0) := (others => '0');
signal s918 : std_logic_vector(33 downto 0) := (others => '0');
signal s919 : std_logic_vector(33 downto 0) := (others => '0');
signal s920 : std_logic_vector(33 downto 0) := (others => '0');
signal s921 : std_logic_vector(33 downto 0) := (others => '0');
signal s922 : std_logic_vector(33 downto 0) := (others => '0');
signal s923 : std_logic_vector(33 downto 0) := (others => '0');
signal s924 : std_logic_vector(33 downto 0) := (others => '0');
signal s925 : std_logic_vector(33 downto 0) := (others => '0');
signal s926 : std_logic_vector(33 downto 0) := (others => '0');
signal s927 : std_logic_vector(33 downto 0) := (others => '0');
signal s928 : std_logic_vector(33 downto 0) := (others => '0');
signal s929 : std_logic_vector(33 downto 0) := (others => '0');
signal s930 : std_logic_vector(33 downto 0) := (others => '0');
signal s931 : std_logic_vector(33 downto 0) := (others => '0');
signal s932 : std_logic_vector(33 downto 0) := (others => '0');
signal s933 : std_logic_vector(33 downto 0) := (others => '0');
signal s934 : std_logic_vector(33 downto 0) := (others => '0');
signal s935 : std_logic_vector(33 downto 0) := (others => '0');
signal s936 : std_logic_vector(33 downto 0) := (others => '0');
signal s937 : std_logic_vector(33 downto 0) := (others => '0');
signal s938 : std_logic_vector(33 downto 0) := (others => '0');
signal s939 : std_logic_vector(33 downto 0) := (others => '0');
signal s940 : std_logic_vector(33 downto 0) := (others => '0');
signal s941 : std_logic_vector(33 downto 0) := (others => '0');
signal s942 : std_logic_vector(33 downto 0) := (others => '0');
signal s943 : std_logic_vector(33 downto 0) := (others => '0');
signal s944 : std_logic_vector(33 downto 0) := (others => '0');
signal s945 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
      s558 <= "0000000000000000000000000000000000";
      s559 <= "0000000000000000000000000000000000";
      s560 <= "0000000000000000000000000000000000";
      s561 <= "0000000000000000000000000000000000";
      s562 <= "0000000000000000000000000000000000";
      s563 <= "0000000000000000000000000000000000";
      s564 <= "0000000000000000000000000000000000";
      s565 <= "0000000000000000000000000000000000";
      s566 <= "0000000000000000000000000000000000";
      s567 <= "0000000000000000000000000000000000";
      s568 <= "0000000000000000000000000000000000";
      s569 <= "0000000000000000000000000000000000";
      s570 <= "0000000000000000000000000000000000";
      s571 <= "0000000000000000000000000000000000";
      s572 <= "0000000000000000000000000000000000";
      s573 <= "0000000000000000000000000000000000";
      s574 <= "0000000000000000000000000000000000";
      s575 <= "0000000000000000000000000000000000";
      s576 <= "0000000000000000000000000000000000";
      s577 <= "0000000000000000000000000000000000";
      s578 <= "0000000000000000000000000000000000";
      s579 <= "0000000000000000000000000000000000";
      s580 <= "0000000000000000000000000000000000";
      s581 <= "0000000000000000000000000000000000";
      s582 <= "0000000000000000000000000000000000";
      s583 <= "0000000000000000000000000000000000";
      s584 <= "0000000000000000000000000000000000";
      s585 <= "0000000000000000000000000000000000";
      s586 <= "0000000000000000000000000000000000";
      s587 <= "0000000000000000000000000000000000";
      s588 <= "0000000000000000000000000000000000";
      s589 <= "0000000000000000000000000000000000";
      s590 <= "0000000000000000000000000000000000";
      s591 <= "0000000000000000000000000000000000";
      s592 <= "0000000000000000000000000000000000";
      s593 <= "0000000000000000000000000000000000";
      s594 <= "0000000000000000000000000000000000";
      s595 <= "0000000000000000000000000000000000";
      s596 <= "0000000000000000000000000000000000";
      s597 <= "0000000000000000000000000000000000";
      s598 <= "0000000000000000000000000000000000";
      s599 <= "0000000000000000000000000000000000";
      s600 <= "0000000000000000000000000000000000";
      s601 <= "0000000000000000000000000000000000";
      s602 <= "0000000000000000000000000000000000";
      s603 <= "0000000000000000000000000000000000";
      s604 <= "0000000000000000000000000000000000";
      s605 <= "0000000000000000000000000000000000";
      s606 <= "0000000000000000000000000000000000";
      s607 <= "0000000000000000000000000000000000";
      s608 <= "0000000000000000000000000000000000";
      s609 <= "0000000000000000000000000000000000";
      s610 <= "0000000000000000000000000000000000";
      s611 <= "0000000000000000000000000000000000";
      s612 <= "0000000000000000000000000000000000";
      s613 <= "0000000000000000000000000000000000";
      s614 <= "0000000000000000000000000000000000";
      s615 <= "0000000000000000000000000000000000";
      s616 <= "0000000000000000000000000000000000";
      s617 <= "0000000000000000000000000000000000";
      s618 <= "0000000000000000000000000000000000";
      s619 <= "0000000000000000000000000000000000";
      s620 <= "0000000000000000000000000000000000";
      s621 <= "0000000000000000000000000000000000";
      s622 <= "0000000000000000000000000000000000";
      s623 <= "0000000000000000000000000000000000";
      s624 <= "0000000000000000000000000000000000";
      s625 <= "0000000000000000000000000000000000";
      s626 <= "0000000000000000000000000000000000";
      s627 <= "0000000000000000000000000000000000";
      s628 <= "0000000000000000000000000000000000";
      s629 <= "0000000000000000000000000000000000";
      s630 <= "0000000000000000000000000000000000";
      s631 <= "0000000000000000000000000000000000";
      s632 <= "0000000000000000000000000000000000";
      s633 <= "0000000000000000000000000000000000";
      s634 <= "0000000000000000000000000000000000";
      s635 <= "0000000000000000000000000000000000";
      s636 <= "0000000000000000000000000000000000";
      s637 <= "0000000000000000000000000000000000";
      s638 <= "0000000000000000000000000000000000";
      s639 <= "0000000000000000000000000000000000";
      s640 <= "0000000000000000000000000000000000";
      s641 <= "0000000000000000000000000000000000";
      s642 <= "0000000000000000000000000000000000";
      s643 <= "0000000000000000000000000000000000";
      s644 <= "0000000000000000000000000000000000";
      s645 <= "0000000000000000000000000000000000";
      s646 <= "0000000000000000000000000000000000";
      s647 <= "0000000000000000000000000000000000";
      s648 <= "0000000000000000000000000000000000";
      s649 <= "0000000000000000000000000000000000";
      s650 <= "0000000000000000000000000000000000";
      s651 <= "0000000000000000000000000000000000";
      s652 <= "0000000000000000000000000000000000";
      s653 <= "0000000000000000000000000000000000";
      s654 <= "0000000000000000000000000000000000";
      s655 <= "0000000000000000000000000000000000";
      s656 <= "0000000000000000000000000000000000";
      s657 <= "0000000000000000000000000000000000";
      s658 <= "0000000000000000000000000000000000";
      s659 <= "0000000000000000000000000000000000";
      s660 <= "0000000000000000000000000000000000";
      s661 <= "0000000000000000000000000000000000";
      s662 <= "0000000000000000000000000000000000";
      s663 <= "0000000000000000000000000000000000";
      s664 <= "0000000000000000000000000000000000";
      s665 <= "0000000000000000000000000000000000";
      s666 <= "0000000000000000000000000000000000";
      s667 <= "0000000000000000000000000000000000";
      s668 <= "0000000000000000000000000000000000";
      s669 <= "0000000000000000000000000000000000";
      s670 <= "0000000000000000000000000000000000";
      s671 <= "0000000000000000000000000000000000";
      s672 <= "0000000000000000000000000000000000";
      s673 <= "0000000000000000000000000000000000";
      s674 <= "0000000000000000000000000000000000";
      s675 <= "0000000000000000000000000000000000";
      s676 <= "0000000000000000000000000000000000";
      s677 <= "0000000000000000000000000000000000";
      s678 <= "0000000000000000000000000000000000";
      s679 <= "0000000000000000000000000000000000";
      s680 <= "0000000000000000000000000000000000";
      s681 <= "0000000000000000000000000000000000";
      s682 <= "0000000000000000000000000000000000";
      s683 <= "0000000000000000000000000000000000";
      s684 <= "0000000000000000000000000000000000";
      s685 <= "0000000000000000000000000000000000";
      s686 <= "0000000000000000000000000000000000";
      s687 <= "0000000000000000000000000000000000";
      s688 <= "0000000000000000000000000000000000";
      s689 <= "0000000000000000000000000000000000";
      s690 <= "0000000000000000000000000000000000";
      s691 <= "0000000000000000000000000000000000";
      s692 <= "0000000000000000000000000000000000";
      s693 <= "0000000000000000000000000000000000";
      s694 <= "0000000000000000000000000000000000";
      s695 <= "0000000000000000000000000000000000";
      s696 <= "0000000000000000000000000000000000";
      s697 <= "0000000000000000000000000000000000";
      s698 <= "0000000000000000000000000000000000";
      s699 <= "0000000000000000000000000000000000";
      s700 <= "0000000000000000000000000000000000";
      s701 <= "0000000000000000000000000000000000";
      s702 <= "0000000000000000000000000000000000";
      s703 <= "0000000000000000000000000000000000";
      s704 <= "0000000000000000000000000000000000";
      s705 <= "0000000000000000000000000000000000";
      s706 <= "0000000000000000000000000000000000";
      s707 <= "0000000000000000000000000000000000";
      s708 <= "0000000000000000000000000000000000";
      s709 <= "0000000000000000000000000000000000";
      s710 <= "0000000000000000000000000000000000";
      s711 <= "0000000000000000000000000000000000";
      s712 <= "0000000000000000000000000000000000";
      s713 <= "0000000000000000000000000000000000";
      s714 <= "0000000000000000000000000000000000";
      s715 <= "0000000000000000000000000000000000";
      s716 <= "0000000000000000000000000000000000";
      s717 <= "0000000000000000000000000000000000";
      s718 <= "0000000000000000000000000000000000";
      s719 <= "0000000000000000000000000000000000";
      s720 <= "0000000000000000000000000000000000";
      s721 <= "0000000000000000000000000000000000";
      s722 <= "0000000000000000000000000000000000";
      s723 <= "0000000000000000000000000000000000";
      s724 <= "0000000000000000000000000000000000";
      s725 <= "0000000000000000000000000000000000";
      s726 <= "0000000000000000000000000000000000";
      s727 <= "0000000000000000000000000000000000";
      s728 <= "0000000000000000000000000000000000";
      s729 <= "0000000000000000000000000000000000";
      s730 <= "0000000000000000000000000000000000";
      s731 <= "0000000000000000000000000000000000";
      s732 <= "0000000000000000000000000000000000";
      s733 <= "0000000000000000000000000000000000";
      s734 <= "0000000000000000000000000000000000";
      s735 <= "0000000000000000000000000000000000";
      s736 <= "0000000000000000000000000000000000";
      s737 <= "0000000000000000000000000000000000";
      s738 <= "0000000000000000000000000000000000";
      s739 <= "0000000000000000000000000000000000";
      s740 <= "0000000000000000000000000000000000";
      s741 <= "0000000000000000000000000000000000";
      s742 <= "0000000000000000000000000000000000";
      s743 <= "0000000000000000000000000000000000";
      s744 <= "0000000000000000000000000000000000";
      s745 <= "0000000000000000000000000000000000";
      s746 <= "0000000000000000000000000000000000";
      s747 <= "0000000000000000000000000000000000";
      s748 <= "0000000000000000000000000000000000";
      s749 <= "0000000000000000000000000000000000";
      s750 <= "0000000000000000000000000000000000";
      s751 <= "0000000000000000000000000000000000";
      s752 <= "0000000000000000000000000000000000";
      s753 <= "0000000000000000000000000000000000";
      s754 <= "0000000000000000000000000000000000";
      s755 <= "0000000000000000000000000000000000";
      s756 <= "0000000000000000000000000000000000";
      s757 <= "0000000000000000000000000000000000";
      s758 <= "0000000000000000000000000000000000";
      s759 <= "0000000000000000000000000000000000";
      s760 <= "0000000000000000000000000000000000";
      s761 <= "0000000000000000000000000000000000";
      s762 <= "0000000000000000000000000000000000";
      s763 <= "0000000000000000000000000000000000";
      s764 <= "0000000000000000000000000000000000";
      s765 <= "0000000000000000000000000000000000";
      s766 <= "0000000000000000000000000000000000";
      s767 <= "0000000000000000000000000000000000";
      s768 <= "0000000000000000000000000000000000";
      s769 <= "0000000000000000000000000000000000";
      s770 <= "0000000000000000000000000000000000";
      s771 <= "0000000000000000000000000000000000";
      s772 <= "0000000000000000000000000000000000";
      s773 <= "0000000000000000000000000000000000";
      s774 <= "0000000000000000000000000000000000";
      s775 <= "0000000000000000000000000000000000";
      s776 <= "0000000000000000000000000000000000";
      s777 <= "0000000000000000000000000000000000";
      s778 <= "0000000000000000000000000000000000";
      s779 <= "0000000000000000000000000000000000";
      s780 <= "0000000000000000000000000000000000";
      s781 <= "0000000000000000000000000000000000";
      s782 <= "0000000000000000000000000000000000";
      s783 <= "0000000000000000000000000000000000";
      s784 <= "0000000000000000000000000000000000";
      s785 <= "0000000000000000000000000000000000";
      s786 <= "0000000000000000000000000000000000";
      s787 <= "0000000000000000000000000000000000";
      s788 <= "0000000000000000000000000000000000";
      s789 <= "0000000000000000000000000000000000";
      s790 <= "0000000000000000000000000000000000";
      s791 <= "0000000000000000000000000000000000";
      s792 <= "0000000000000000000000000000000000";
      s793 <= "0000000000000000000000000000000000";
      s794 <= "0000000000000000000000000000000000";
      s795 <= "0000000000000000000000000000000000";
      s796 <= "0000000000000000000000000000000000";
      s797 <= "0000000000000000000000000000000000";
      s798 <= "0000000000000000000000000000000000";
      s799 <= "0000000000000000000000000000000000";
      s800 <= "0000000000000000000000000000000000";
      s801 <= "0000000000000000000000000000000000";
      s802 <= "0000000000000000000000000000000000";
      s803 <= "0000000000000000000000000000000000";
      s804 <= "0000000000000000000000000000000000";
      s805 <= "0000000000000000000000000000000000";
      s806 <= "0000000000000000000000000000000000";
      s807 <= "0000000000000000000000000000000000";
      s808 <= "0000000000000000000000000000000000";
      s809 <= "0000000000000000000000000000000000";
      s810 <= "0000000000000000000000000000000000";
      s811 <= "0000000000000000000000000000000000";
      s812 <= "0000000000000000000000000000000000";
      s813 <= "0000000000000000000000000000000000";
      s814 <= "0000000000000000000000000000000000";
      s815 <= "0000000000000000000000000000000000";
      s816 <= "0000000000000000000000000000000000";
      s817 <= "0000000000000000000000000000000000";
      s818 <= "0000000000000000000000000000000000";
      s819 <= "0000000000000000000000000000000000";
      s820 <= "0000000000000000000000000000000000";
      s821 <= "0000000000000000000000000000000000";
      s822 <= "0000000000000000000000000000000000";
      s823 <= "0000000000000000000000000000000000";
      s824 <= "0000000000000000000000000000000000";
      s825 <= "0000000000000000000000000000000000";
      s826 <= "0000000000000000000000000000000000";
      s827 <= "0000000000000000000000000000000000";
      s828 <= "0000000000000000000000000000000000";
      s829 <= "0000000000000000000000000000000000";
      s830 <= "0000000000000000000000000000000000";
      s831 <= "0000000000000000000000000000000000";
      s832 <= "0000000000000000000000000000000000";
      s833 <= "0000000000000000000000000000000000";
      s834 <= "0000000000000000000000000000000000";
      s835 <= "0000000000000000000000000000000000";
      s836 <= "0000000000000000000000000000000000";
      s837 <= "0000000000000000000000000000000000";
      s838 <= "0000000000000000000000000000000000";
      s839 <= "0000000000000000000000000000000000";
      s840 <= "0000000000000000000000000000000000";
      s841 <= "0000000000000000000000000000000000";
      s842 <= "0000000000000000000000000000000000";
      s843 <= "0000000000000000000000000000000000";
      s844 <= "0000000000000000000000000000000000";
      s845 <= "0000000000000000000000000000000000";
      s846 <= "0000000000000000000000000000000000";
      s847 <= "0000000000000000000000000000000000";
      s848 <= "0000000000000000000000000000000000";
      s849 <= "0000000000000000000000000000000000";
      s850 <= "0000000000000000000000000000000000";
      s851 <= "0000000000000000000000000000000000";
      s852 <= "0000000000000000000000000000000000";
      s853 <= "0000000000000000000000000000000000";
      s854 <= "0000000000000000000000000000000000";
      s855 <= "0000000000000000000000000000000000";
      s856 <= "0000000000000000000000000000000000";
      s857 <= "0000000000000000000000000000000000";
      s858 <= "0000000000000000000000000000000000";
      s859 <= "0000000000000000000000000000000000";
      s860 <= "0000000000000000000000000000000000";
      s861 <= "0000000000000000000000000000000000";
      s862 <= "0000000000000000000000000000000000";
      s863 <= "0000000000000000000000000000000000";
      s864 <= "0000000000000000000000000000000000";
      s865 <= "0000000000000000000000000000000000";
      s866 <= "0000000000000000000000000000000000";
      s867 <= "0000000000000000000000000000000000";
      s868 <= "0000000000000000000000000000000000";
      s869 <= "0000000000000000000000000000000000";
      s870 <= "0000000000000000000000000000000000";
      s871 <= "0000000000000000000000000000000000";
      s872 <= "0000000000000000000000000000000000";
      s873 <= "0000000000000000000000000000000000";
      s874 <= "0000000000000000000000000000000000";
      s875 <= "0000000000000000000000000000000000";
      s876 <= "0000000000000000000000000000000000";
      s877 <= "0000000000000000000000000000000000";
      s878 <= "0000000000000000000000000000000000";
      s879 <= "0000000000000000000000000000000000";
      s880 <= "0000000000000000000000000000000000";
      s881 <= "0000000000000000000000000000000000";
      s882 <= "0000000000000000000000000000000000";
      s883 <= "0000000000000000000000000000000000";
      s884 <= "0000000000000000000000000000000000";
      s885 <= "0000000000000000000000000000000000";
      s886 <= "0000000000000000000000000000000000";
      s887 <= "0000000000000000000000000000000000";
      s888 <= "0000000000000000000000000000000000";
      s889 <= "0000000000000000000000000000000000";
      s890 <= "0000000000000000000000000000000000";
      s891 <= "0000000000000000000000000000000000";
      s892 <= "0000000000000000000000000000000000";
      s893 <= "0000000000000000000000000000000000";
      s894 <= "0000000000000000000000000000000000";
      s895 <= "0000000000000000000000000000000000";
      s896 <= "0000000000000000000000000000000000";
      s897 <= "0000000000000000000000000000000000";
      s898 <= "0000000000000000000000000000000000";
      s899 <= "0000000000000000000000000000000000";
      s900 <= "0000000000000000000000000000000000";
      s901 <= "0000000000000000000000000000000000";
      s902 <= "0000000000000000000000000000000000";
      s903 <= "0000000000000000000000000000000000";
      s904 <= "0000000000000000000000000000000000";
      s905 <= "0000000000000000000000000000000000";
      s906 <= "0000000000000000000000000000000000";
      s907 <= "0000000000000000000000000000000000";
      s908 <= "0000000000000000000000000000000000";
      s909 <= "0000000000000000000000000000000000";
      s910 <= "0000000000000000000000000000000000";
      s911 <= "0000000000000000000000000000000000";
      s912 <= "0000000000000000000000000000000000";
      s913 <= "0000000000000000000000000000000000";
      s914 <= "0000000000000000000000000000000000";
      s915 <= "0000000000000000000000000000000000";
      s916 <= "0000000000000000000000000000000000";
      s917 <= "0000000000000000000000000000000000";
      s918 <= "0000000000000000000000000000000000";
      s919 <= "0000000000000000000000000000000000";
      s920 <= "0000000000000000000000000000000000";
      s921 <= "0000000000000000000000000000000000";
      s922 <= "0000000000000000000000000000000000";
      s923 <= "0000000000000000000000000000000000";
      s924 <= "0000000000000000000000000000000000";
      s925 <= "0000000000000000000000000000000000";
      s926 <= "0000000000000000000000000000000000";
      s927 <= "0000000000000000000000000000000000";
      s928 <= "0000000000000000000000000000000000";
      s929 <= "0000000000000000000000000000000000";
      s930 <= "0000000000000000000000000000000000";
      s931 <= "0000000000000000000000000000000000";
      s932 <= "0000000000000000000000000000000000";
      s933 <= "0000000000000000000000000000000000";
      s934 <= "0000000000000000000000000000000000";
      s935 <= "0000000000000000000000000000000000";
      s936 <= "0000000000000000000000000000000000";
      s937 <= "0000000000000000000000000000000000";
      s938 <= "0000000000000000000000000000000000";
      s939 <= "0000000000000000000000000000000000";
      s940 <= "0000000000000000000000000000000000";
      s941 <= "0000000000000000000000000000000000";
      s942 <= "0000000000000000000000000000000000";
      s943 <= "0000000000000000000000000000000000";
      s944 <= "0000000000000000000000000000000000";
      s945 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      s558 <= s557;
      s559 <= s558;
      s560 <= s559;
      s561 <= s560;
      s562 <= s561;
      s563 <= s562;
      s564 <= s563;
      s565 <= s564;
      s566 <= s565;
      s567 <= s566;
      s568 <= s567;
      s569 <= s568;
      s570 <= s569;
      s571 <= s570;
      s572 <= s571;
      s573 <= s572;
      s574 <= s573;
      s575 <= s574;
      s576 <= s575;
      s577 <= s576;
      s578 <= s577;
      s579 <= s578;
      s580 <= s579;
      s581 <= s580;
      s582 <= s581;
      s583 <= s582;
      s584 <= s583;
      s585 <= s584;
      s586 <= s585;
      s587 <= s586;
      s588 <= s587;
      s589 <= s588;
      s590 <= s589;
      s591 <= s590;
      s592 <= s591;
      s593 <= s592;
      s594 <= s593;
      s595 <= s594;
      s596 <= s595;
      s597 <= s596;
      s598 <= s597;
      s599 <= s598;
      s600 <= s599;
      s601 <= s600;
      s602 <= s601;
      s603 <= s602;
      s604 <= s603;
      s605 <= s604;
      s606 <= s605;
      s607 <= s606;
      s608 <= s607;
      s609 <= s608;
      s610 <= s609;
      s611 <= s610;
      s612 <= s611;
      s613 <= s612;
      s614 <= s613;
      s615 <= s614;
      s616 <= s615;
      s617 <= s616;
      s618 <= s617;
      s619 <= s618;
      s620 <= s619;
      s621 <= s620;
      s622 <= s621;
      s623 <= s622;
      s624 <= s623;
      s625 <= s624;
      s626 <= s625;
      s627 <= s626;
      s628 <= s627;
      s629 <= s628;
      s630 <= s629;
      s631 <= s630;
      s632 <= s631;
      s633 <= s632;
      s634 <= s633;
      s635 <= s634;
      s636 <= s635;
      s637 <= s636;
      s638 <= s637;
      s639 <= s638;
      s640 <= s639;
      s641 <= s640;
      s642 <= s641;
      s643 <= s642;
      s644 <= s643;
      s645 <= s644;
      s646 <= s645;
      s647 <= s646;
      s648 <= s647;
      s649 <= s648;
      s650 <= s649;
      s651 <= s650;
      s652 <= s651;
      s653 <= s652;
      s654 <= s653;
      s655 <= s654;
      s656 <= s655;
      s657 <= s656;
      s658 <= s657;
      s659 <= s658;
      s660 <= s659;
      s661 <= s660;
      s662 <= s661;
      s663 <= s662;
      s664 <= s663;
      s665 <= s664;
      s666 <= s665;
      s667 <= s666;
      s668 <= s667;
      s669 <= s668;
      s670 <= s669;
      s671 <= s670;
      s672 <= s671;
      s673 <= s672;
      s674 <= s673;
      s675 <= s674;
      s676 <= s675;
      s677 <= s676;
      s678 <= s677;
      s679 <= s678;
      s680 <= s679;
      s681 <= s680;
      s682 <= s681;
      s683 <= s682;
      s684 <= s683;
      s685 <= s684;
      s686 <= s685;
      s687 <= s686;
      s688 <= s687;
      s689 <= s688;
      s690 <= s689;
      s691 <= s690;
      s692 <= s691;
      s693 <= s692;
      s694 <= s693;
      s695 <= s694;
      s696 <= s695;
      s697 <= s696;
      s698 <= s697;
      s699 <= s698;
      s700 <= s699;
      s701 <= s700;
      s702 <= s701;
      s703 <= s702;
      s704 <= s703;
      s705 <= s704;
      s706 <= s705;
      s707 <= s706;
      s708 <= s707;
      s709 <= s708;
      s710 <= s709;
      s711 <= s710;
      s712 <= s711;
      s713 <= s712;
      s714 <= s713;
      s715 <= s714;
      s716 <= s715;
      s717 <= s716;
      s718 <= s717;
      s719 <= s718;
      s720 <= s719;
      s721 <= s720;
      s722 <= s721;
      s723 <= s722;
      s724 <= s723;
      s725 <= s724;
      s726 <= s725;
      s727 <= s726;
      s728 <= s727;
      s729 <= s728;
      s730 <= s729;
      s731 <= s730;
      s732 <= s731;
      s733 <= s732;
      s734 <= s733;
      s735 <= s734;
      s736 <= s735;
      s737 <= s736;
      s738 <= s737;
      s739 <= s738;
      s740 <= s739;
      s741 <= s740;
      s742 <= s741;
      s743 <= s742;
      s744 <= s743;
      s745 <= s744;
      s746 <= s745;
      s747 <= s746;
      s748 <= s747;
      s749 <= s748;
      s750 <= s749;
      s751 <= s750;
      s752 <= s751;
      s753 <= s752;
      s754 <= s753;
      s755 <= s754;
      s756 <= s755;
      s757 <= s756;
      s758 <= s757;
      s759 <= s758;
      s760 <= s759;
      s761 <= s760;
      s762 <= s761;
      s763 <= s762;
      s764 <= s763;
      s765 <= s764;
      s766 <= s765;
      s767 <= s766;
      s768 <= s767;
      s769 <= s768;
      s770 <= s769;
      s771 <= s770;
      s772 <= s771;
      s773 <= s772;
      s774 <= s773;
      s775 <= s774;
      s776 <= s775;
      s777 <= s776;
      s778 <= s777;
      s779 <= s778;
      s780 <= s779;
      s781 <= s780;
      s782 <= s781;
      s783 <= s782;
      s784 <= s783;
      s785 <= s784;
      s786 <= s785;
      s787 <= s786;
      s788 <= s787;
      s789 <= s788;
      s790 <= s789;
      s791 <= s790;
      s792 <= s791;
      s793 <= s792;
      s794 <= s793;
      s795 <= s794;
      s796 <= s795;
      s797 <= s796;
      s798 <= s797;
      s799 <= s798;
      s800 <= s799;
      s801 <= s800;
      s802 <= s801;
      s803 <= s802;
      s804 <= s803;
      s805 <= s804;
      s806 <= s805;
      s807 <= s806;
      s808 <= s807;
      s809 <= s808;
      s810 <= s809;
      s811 <= s810;
      s812 <= s811;
      s813 <= s812;
      s814 <= s813;
      s815 <= s814;
      s816 <= s815;
      s817 <= s816;
      s818 <= s817;
      s819 <= s818;
      s820 <= s819;
      s821 <= s820;
      s822 <= s821;
      s823 <= s822;
      s824 <= s823;
      s825 <= s824;
      s826 <= s825;
      s827 <= s826;
      s828 <= s827;
      s829 <= s828;
      s830 <= s829;
      s831 <= s830;
      s832 <= s831;
      s833 <= s832;
      s834 <= s833;
      s835 <= s834;
      s836 <= s835;
      s837 <= s836;
      s838 <= s837;
      s839 <= s838;
      s840 <= s839;
      s841 <= s840;
      s842 <= s841;
      s843 <= s842;
      s844 <= s843;
      s845 <= s844;
      s846 <= s845;
      s847 <= s846;
      s848 <= s847;
      s849 <= s848;
      s850 <= s849;
      s851 <= s850;
      s852 <= s851;
      s853 <= s852;
      s854 <= s853;
      s855 <= s854;
      s856 <= s855;
      s857 <= s856;
      s858 <= s857;
      s859 <= s858;
      s860 <= s859;
      s861 <= s860;
      s862 <= s861;
      s863 <= s862;
      s864 <= s863;
      s865 <= s864;
      s866 <= s865;
      s867 <= s866;
      s868 <= s867;
      s869 <= s868;
      s870 <= s869;
      s871 <= s870;
      s872 <= s871;
      s873 <= s872;
      s874 <= s873;
      s875 <= s874;
      s876 <= s875;
      s877 <= s876;
      s878 <= s877;
      s879 <= s878;
      s880 <= s879;
      s881 <= s880;
      s882 <= s881;
      s883 <= s882;
      s884 <= s883;
      s885 <= s884;
      s886 <= s885;
      s887 <= s886;
      s888 <= s887;
      s889 <= s888;
      s890 <= s889;
      s891 <= s890;
      s892 <= s891;
      s893 <= s892;
      s894 <= s893;
      s895 <= s894;
      s896 <= s895;
      s897 <= s896;
      s898 <= s897;
      s899 <= s898;
      s900 <= s899;
      s901 <= s900;
      s902 <= s901;
      s903 <= s902;
      s904 <= s903;
      s905 <= s904;
      s906 <= s905;
      s907 <= s906;
      s908 <= s907;
      s909 <= s908;
      s910 <= s909;
      s911 <= s910;
      s912 <= s911;
      s913 <= s912;
      s914 <= s913;
      s915 <= s914;
      s916 <= s915;
      s917 <= s916;
      s918 <= s917;
      s919 <= s918;
      s920 <= s919;
      s921 <= s920;
      s922 <= s921;
      s923 <= s922;
      s924 <= s923;
      s925 <= s924;
      s926 <= s925;
      s927 <= s926;
      s928 <= s927;
      s929 <= s928;
      s930 <= s929;
      s931 <= s930;
      s932 <= s931;
      s933 <= s932;
      s934 <= s933;
      s935 <= s934;
      s936 <= s935;
      s937 <= s936;
      s938 <= s937;
      s939 <= s938;
      s940 <= s939;
      s941 <= s940;
      s942 <= s941;
      s943 <= s942;
      s944 <= s943;
      s945 <= s944;
      Y <= s945;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_995_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 995 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_995_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_995_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
signal s558 : std_logic_vector(33 downto 0) := (others => '0');
signal s559 : std_logic_vector(33 downto 0) := (others => '0');
signal s560 : std_logic_vector(33 downto 0) := (others => '0');
signal s561 : std_logic_vector(33 downto 0) := (others => '0');
signal s562 : std_logic_vector(33 downto 0) := (others => '0');
signal s563 : std_logic_vector(33 downto 0) := (others => '0');
signal s564 : std_logic_vector(33 downto 0) := (others => '0');
signal s565 : std_logic_vector(33 downto 0) := (others => '0');
signal s566 : std_logic_vector(33 downto 0) := (others => '0');
signal s567 : std_logic_vector(33 downto 0) := (others => '0');
signal s568 : std_logic_vector(33 downto 0) := (others => '0');
signal s569 : std_logic_vector(33 downto 0) := (others => '0');
signal s570 : std_logic_vector(33 downto 0) := (others => '0');
signal s571 : std_logic_vector(33 downto 0) := (others => '0');
signal s572 : std_logic_vector(33 downto 0) := (others => '0');
signal s573 : std_logic_vector(33 downto 0) := (others => '0');
signal s574 : std_logic_vector(33 downto 0) := (others => '0');
signal s575 : std_logic_vector(33 downto 0) := (others => '0');
signal s576 : std_logic_vector(33 downto 0) := (others => '0');
signal s577 : std_logic_vector(33 downto 0) := (others => '0');
signal s578 : std_logic_vector(33 downto 0) := (others => '0');
signal s579 : std_logic_vector(33 downto 0) := (others => '0');
signal s580 : std_logic_vector(33 downto 0) := (others => '0');
signal s581 : std_logic_vector(33 downto 0) := (others => '0');
signal s582 : std_logic_vector(33 downto 0) := (others => '0');
signal s583 : std_logic_vector(33 downto 0) := (others => '0');
signal s584 : std_logic_vector(33 downto 0) := (others => '0');
signal s585 : std_logic_vector(33 downto 0) := (others => '0');
signal s586 : std_logic_vector(33 downto 0) := (others => '0');
signal s587 : std_logic_vector(33 downto 0) := (others => '0');
signal s588 : std_logic_vector(33 downto 0) := (others => '0');
signal s589 : std_logic_vector(33 downto 0) := (others => '0');
signal s590 : std_logic_vector(33 downto 0) := (others => '0');
signal s591 : std_logic_vector(33 downto 0) := (others => '0');
signal s592 : std_logic_vector(33 downto 0) := (others => '0');
signal s593 : std_logic_vector(33 downto 0) := (others => '0');
signal s594 : std_logic_vector(33 downto 0) := (others => '0');
signal s595 : std_logic_vector(33 downto 0) := (others => '0');
signal s596 : std_logic_vector(33 downto 0) := (others => '0');
signal s597 : std_logic_vector(33 downto 0) := (others => '0');
signal s598 : std_logic_vector(33 downto 0) := (others => '0');
signal s599 : std_logic_vector(33 downto 0) := (others => '0');
signal s600 : std_logic_vector(33 downto 0) := (others => '0');
signal s601 : std_logic_vector(33 downto 0) := (others => '0');
signal s602 : std_logic_vector(33 downto 0) := (others => '0');
signal s603 : std_logic_vector(33 downto 0) := (others => '0');
signal s604 : std_logic_vector(33 downto 0) := (others => '0');
signal s605 : std_logic_vector(33 downto 0) := (others => '0');
signal s606 : std_logic_vector(33 downto 0) := (others => '0');
signal s607 : std_logic_vector(33 downto 0) := (others => '0');
signal s608 : std_logic_vector(33 downto 0) := (others => '0');
signal s609 : std_logic_vector(33 downto 0) := (others => '0');
signal s610 : std_logic_vector(33 downto 0) := (others => '0');
signal s611 : std_logic_vector(33 downto 0) := (others => '0');
signal s612 : std_logic_vector(33 downto 0) := (others => '0');
signal s613 : std_logic_vector(33 downto 0) := (others => '0');
signal s614 : std_logic_vector(33 downto 0) := (others => '0');
signal s615 : std_logic_vector(33 downto 0) := (others => '0');
signal s616 : std_logic_vector(33 downto 0) := (others => '0');
signal s617 : std_logic_vector(33 downto 0) := (others => '0');
signal s618 : std_logic_vector(33 downto 0) := (others => '0');
signal s619 : std_logic_vector(33 downto 0) := (others => '0');
signal s620 : std_logic_vector(33 downto 0) := (others => '0');
signal s621 : std_logic_vector(33 downto 0) := (others => '0');
signal s622 : std_logic_vector(33 downto 0) := (others => '0');
signal s623 : std_logic_vector(33 downto 0) := (others => '0');
signal s624 : std_logic_vector(33 downto 0) := (others => '0');
signal s625 : std_logic_vector(33 downto 0) := (others => '0');
signal s626 : std_logic_vector(33 downto 0) := (others => '0');
signal s627 : std_logic_vector(33 downto 0) := (others => '0');
signal s628 : std_logic_vector(33 downto 0) := (others => '0');
signal s629 : std_logic_vector(33 downto 0) := (others => '0');
signal s630 : std_logic_vector(33 downto 0) := (others => '0');
signal s631 : std_logic_vector(33 downto 0) := (others => '0');
signal s632 : std_logic_vector(33 downto 0) := (others => '0');
signal s633 : std_logic_vector(33 downto 0) := (others => '0');
signal s634 : std_logic_vector(33 downto 0) := (others => '0');
signal s635 : std_logic_vector(33 downto 0) := (others => '0');
signal s636 : std_logic_vector(33 downto 0) := (others => '0');
signal s637 : std_logic_vector(33 downto 0) := (others => '0');
signal s638 : std_logic_vector(33 downto 0) := (others => '0');
signal s639 : std_logic_vector(33 downto 0) := (others => '0');
signal s640 : std_logic_vector(33 downto 0) := (others => '0');
signal s641 : std_logic_vector(33 downto 0) := (others => '0');
signal s642 : std_logic_vector(33 downto 0) := (others => '0');
signal s643 : std_logic_vector(33 downto 0) := (others => '0');
signal s644 : std_logic_vector(33 downto 0) := (others => '0');
signal s645 : std_logic_vector(33 downto 0) := (others => '0');
signal s646 : std_logic_vector(33 downto 0) := (others => '0');
signal s647 : std_logic_vector(33 downto 0) := (others => '0');
signal s648 : std_logic_vector(33 downto 0) := (others => '0');
signal s649 : std_logic_vector(33 downto 0) := (others => '0');
signal s650 : std_logic_vector(33 downto 0) := (others => '0');
signal s651 : std_logic_vector(33 downto 0) := (others => '0');
signal s652 : std_logic_vector(33 downto 0) := (others => '0');
signal s653 : std_logic_vector(33 downto 0) := (others => '0');
signal s654 : std_logic_vector(33 downto 0) := (others => '0');
signal s655 : std_logic_vector(33 downto 0) := (others => '0');
signal s656 : std_logic_vector(33 downto 0) := (others => '0');
signal s657 : std_logic_vector(33 downto 0) := (others => '0');
signal s658 : std_logic_vector(33 downto 0) := (others => '0');
signal s659 : std_logic_vector(33 downto 0) := (others => '0');
signal s660 : std_logic_vector(33 downto 0) := (others => '0');
signal s661 : std_logic_vector(33 downto 0) := (others => '0');
signal s662 : std_logic_vector(33 downto 0) := (others => '0');
signal s663 : std_logic_vector(33 downto 0) := (others => '0');
signal s664 : std_logic_vector(33 downto 0) := (others => '0');
signal s665 : std_logic_vector(33 downto 0) := (others => '0');
signal s666 : std_logic_vector(33 downto 0) := (others => '0');
signal s667 : std_logic_vector(33 downto 0) := (others => '0');
signal s668 : std_logic_vector(33 downto 0) := (others => '0');
signal s669 : std_logic_vector(33 downto 0) := (others => '0');
signal s670 : std_logic_vector(33 downto 0) := (others => '0');
signal s671 : std_logic_vector(33 downto 0) := (others => '0');
signal s672 : std_logic_vector(33 downto 0) := (others => '0');
signal s673 : std_logic_vector(33 downto 0) := (others => '0');
signal s674 : std_logic_vector(33 downto 0) := (others => '0');
signal s675 : std_logic_vector(33 downto 0) := (others => '0');
signal s676 : std_logic_vector(33 downto 0) := (others => '0');
signal s677 : std_logic_vector(33 downto 0) := (others => '0');
signal s678 : std_logic_vector(33 downto 0) := (others => '0');
signal s679 : std_logic_vector(33 downto 0) := (others => '0');
signal s680 : std_logic_vector(33 downto 0) := (others => '0');
signal s681 : std_logic_vector(33 downto 0) := (others => '0');
signal s682 : std_logic_vector(33 downto 0) := (others => '0');
signal s683 : std_logic_vector(33 downto 0) := (others => '0');
signal s684 : std_logic_vector(33 downto 0) := (others => '0');
signal s685 : std_logic_vector(33 downto 0) := (others => '0');
signal s686 : std_logic_vector(33 downto 0) := (others => '0');
signal s687 : std_logic_vector(33 downto 0) := (others => '0');
signal s688 : std_logic_vector(33 downto 0) := (others => '0');
signal s689 : std_logic_vector(33 downto 0) := (others => '0');
signal s690 : std_logic_vector(33 downto 0) := (others => '0');
signal s691 : std_logic_vector(33 downto 0) := (others => '0');
signal s692 : std_logic_vector(33 downto 0) := (others => '0');
signal s693 : std_logic_vector(33 downto 0) := (others => '0');
signal s694 : std_logic_vector(33 downto 0) := (others => '0');
signal s695 : std_logic_vector(33 downto 0) := (others => '0');
signal s696 : std_logic_vector(33 downto 0) := (others => '0');
signal s697 : std_logic_vector(33 downto 0) := (others => '0');
signal s698 : std_logic_vector(33 downto 0) := (others => '0');
signal s699 : std_logic_vector(33 downto 0) := (others => '0');
signal s700 : std_logic_vector(33 downto 0) := (others => '0');
signal s701 : std_logic_vector(33 downto 0) := (others => '0');
signal s702 : std_logic_vector(33 downto 0) := (others => '0');
signal s703 : std_logic_vector(33 downto 0) := (others => '0');
signal s704 : std_logic_vector(33 downto 0) := (others => '0');
signal s705 : std_logic_vector(33 downto 0) := (others => '0');
signal s706 : std_logic_vector(33 downto 0) := (others => '0');
signal s707 : std_logic_vector(33 downto 0) := (others => '0');
signal s708 : std_logic_vector(33 downto 0) := (others => '0');
signal s709 : std_logic_vector(33 downto 0) := (others => '0');
signal s710 : std_logic_vector(33 downto 0) := (others => '0');
signal s711 : std_logic_vector(33 downto 0) := (others => '0');
signal s712 : std_logic_vector(33 downto 0) := (others => '0');
signal s713 : std_logic_vector(33 downto 0) := (others => '0');
signal s714 : std_logic_vector(33 downto 0) := (others => '0');
signal s715 : std_logic_vector(33 downto 0) := (others => '0');
signal s716 : std_logic_vector(33 downto 0) := (others => '0');
signal s717 : std_logic_vector(33 downto 0) := (others => '0');
signal s718 : std_logic_vector(33 downto 0) := (others => '0');
signal s719 : std_logic_vector(33 downto 0) := (others => '0');
signal s720 : std_logic_vector(33 downto 0) := (others => '0');
signal s721 : std_logic_vector(33 downto 0) := (others => '0');
signal s722 : std_logic_vector(33 downto 0) := (others => '0');
signal s723 : std_logic_vector(33 downto 0) := (others => '0');
signal s724 : std_logic_vector(33 downto 0) := (others => '0');
signal s725 : std_logic_vector(33 downto 0) := (others => '0');
signal s726 : std_logic_vector(33 downto 0) := (others => '0');
signal s727 : std_logic_vector(33 downto 0) := (others => '0');
signal s728 : std_logic_vector(33 downto 0) := (others => '0');
signal s729 : std_logic_vector(33 downto 0) := (others => '0');
signal s730 : std_logic_vector(33 downto 0) := (others => '0');
signal s731 : std_logic_vector(33 downto 0) := (others => '0');
signal s732 : std_logic_vector(33 downto 0) := (others => '0');
signal s733 : std_logic_vector(33 downto 0) := (others => '0');
signal s734 : std_logic_vector(33 downto 0) := (others => '0');
signal s735 : std_logic_vector(33 downto 0) := (others => '0');
signal s736 : std_logic_vector(33 downto 0) := (others => '0');
signal s737 : std_logic_vector(33 downto 0) := (others => '0');
signal s738 : std_logic_vector(33 downto 0) := (others => '0');
signal s739 : std_logic_vector(33 downto 0) := (others => '0');
signal s740 : std_logic_vector(33 downto 0) := (others => '0');
signal s741 : std_logic_vector(33 downto 0) := (others => '0');
signal s742 : std_logic_vector(33 downto 0) := (others => '0');
signal s743 : std_logic_vector(33 downto 0) := (others => '0');
signal s744 : std_logic_vector(33 downto 0) := (others => '0');
signal s745 : std_logic_vector(33 downto 0) := (others => '0');
signal s746 : std_logic_vector(33 downto 0) := (others => '0');
signal s747 : std_logic_vector(33 downto 0) := (others => '0');
signal s748 : std_logic_vector(33 downto 0) := (others => '0');
signal s749 : std_logic_vector(33 downto 0) := (others => '0');
signal s750 : std_logic_vector(33 downto 0) := (others => '0');
signal s751 : std_logic_vector(33 downto 0) := (others => '0');
signal s752 : std_logic_vector(33 downto 0) := (others => '0');
signal s753 : std_logic_vector(33 downto 0) := (others => '0');
signal s754 : std_logic_vector(33 downto 0) := (others => '0');
signal s755 : std_logic_vector(33 downto 0) := (others => '0');
signal s756 : std_logic_vector(33 downto 0) := (others => '0');
signal s757 : std_logic_vector(33 downto 0) := (others => '0');
signal s758 : std_logic_vector(33 downto 0) := (others => '0');
signal s759 : std_logic_vector(33 downto 0) := (others => '0');
signal s760 : std_logic_vector(33 downto 0) := (others => '0');
signal s761 : std_logic_vector(33 downto 0) := (others => '0');
signal s762 : std_logic_vector(33 downto 0) := (others => '0');
signal s763 : std_logic_vector(33 downto 0) := (others => '0');
signal s764 : std_logic_vector(33 downto 0) := (others => '0');
signal s765 : std_logic_vector(33 downto 0) := (others => '0');
signal s766 : std_logic_vector(33 downto 0) := (others => '0');
signal s767 : std_logic_vector(33 downto 0) := (others => '0');
signal s768 : std_logic_vector(33 downto 0) := (others => '0');
signal s769 : std_logic_vector(33 downto 0) := (others => '0');
signal s770 : std_logic_vector(33 downto 0) := (others => '0');
signal s771 : std_logic_vector(33 downto 0) := (others => '0');
signal s772 : std_logic_vector(33 downto 0) := (others => '0');
signal s773 : std_logic_vector(33 downto 0) := (others => '0');
signal s774 : std_logic_vector(33 downto 0) := (others => '0');
signal s775 : std_logic_vector(33 downto 0) := (others => '0');
signal s776 : std_logic_vector(33 downto 0) := (others => '0');
signal s777 : std_logic_vector(33 downto 0) := (others => '0');
signal s778 : std_logic_vector(33 downto 0) := (others => '0');
signal s779 : std_logic_vector(33 downto 0) := (others => '0');
signal s780 : std_logic_vector(33 downto 0) := (others => '0');
signal s781 : std_logic_vector(33 downto 0) := (others => '0');
signal s782 : std_logic_vector(33 downto 0) := (others => '0');
signal s783 : std_logic_vector(33 downto 0) := (others => '0');
signal s784 : std_logic_vector(33 downto 0) := (others => '0');
signal s785 : std_logic_vector(33 downto 0) := (others => '0');
signal s786 : std_logic_vector(33 downto 0) := (others => '0');
signal s787 : std_logic_vector(33 downto 0) := (others => '0');
signal s788 : std_logic_vector(33 downto 0) := (others => '0');
signal s789 : std_logic_vector(33 downto 0) := (others => '0');
signal s790 : std_logic_vector(33 downto 0) := (others => '0');
signal s791 : std_logic_vector(33 downto 0) := (others => '0');
signal s792 : std_logic_vector(33 downto 0) := (others => '0');
signal s793 : std_logic_vector(33 downto 0) := (others => '0');
signal s794 : std_logic_vector(33 downto 0) := (others => '0');
signal s795 : std_logic_vector(33 downto 0) := (others => '0');
signal s796 : std_logic_vector(33 downto 0) := (others => '0');
signal s797 : std_logic_vector(33 downto 0) := (others => '0');
signal s798 : std_logic_vector(33 downto 0) := (others => '0');
signal s799 : std_logic_vector(33 downto 0) := (others => '0');
signal s800 : std_logic_vector(33 downto 0) := (others => '0');
signal s801 : std_logic_vector(33 downto 0) := (others => '0');
signal s802 : std_logic_vector(33 downto 0) := (others => '0');
signal s803 : std_logic_vector(33 downto 0) := (others => '0');
signal s804 : std_logic_vector(33 downto 0) := (others => '0');
signal s805 : std_logic_vector(33 downto 0) := (others => '0');
signal s806 : std_logic_vector(33 downto 0) := (others => '0');
signal s807 : std_logic_vector(33 downto 0) := (others => '0');
signal s808 : std_logic_vector(33 downto 0) := (others => '0');
signal s809 : std_logic_vector(33 downto 0) := (others => '0');
signal s810 : std_logic_vector(33 downto 0) := (others => '0');
signal s811 : std_logic_vector(33 downto 0) := (others => '0');
signal s812 : std_logic_vector(33 downto 0) := (others => '0');
signal s813 : std_logic_vector(33 downto 0) := (others => '0');
signal s814 : std_logic_vector(33 downto 0) := (others => '0');
signal s815 : std_logic_vector(33 downto 0) := (others => '0');
signal s816 : std_logic_vector(33 downto 0) := (others => '0');
signal s817 : std_logic_vector(33 downto 0) := (others => '0');
signal s818 : std_logic_vector(33 downto 0) := (others => '0');
signal s819 : std_logic_vector(33 downto 0) := (others => '0');
signal s820 : std_logic_vector(33 downto 0) := (others => '0');
signal s821 : std_logic_vector(33 downto 0) := (others => '0');
signal s822 : std_logic_vector(33 downto 0) := (others => '0');
signal s823 : std_logic_vector(33 downto 0) := (others => '0');
signal s824 : std_logic_vector(33 downto 0) := (others => '0');
signal s825 : std_logic_vector(33 downto 0) := (others => '0');
signal s826 : std_logic_vector(33 downto 0) := (others => '0');
signal s827 : std_logic_vector(33 downto 0) := (others => '0');
signal s828 : std_logic_vector(33 downto 0) := (others => '0');
signal s829 : std_logic_vector(33 downto 0) := (others => '0');
signal s830 : std_logic_vector(33 downto 0) := (others => '0');
signal s831 : std_logic_vector(33 downto 0) := (others => '0');
signal s832 : std_logic_vector(33 downto 0) := (others => '0');
signal s833 : std_logic_vector(33 downto 0) := (others => '0');
signal s834 : std_logic_vector(33 downto 0) := (others => '0');
signal s835 : std_logic_vector(33 downto 0) := (others => '0');
signal s836 : std_logic_vector(33 downto 0) := (others => '0');
signal s837 : std_logic_vector(33 downto 0) := (others => '0');
signal s838 : std_logic_vector(33 downto 0) := (others => '0');
signal s839 : std_logic_vector(33 downto 0) := (others => '0');
signal s840 : std_logic_vector(33 downto 0) := (others => '0');
signal s841 : std_logic_vector(33 downto 0) := (others => '0');
signal s842 : std_logic_vector(33 downto 0) := (others => '0');
signal s843 : std_logic_vector(33 downto 0) := (others => '0');
signal s844 : std_logic_vector(33 downto 0) := (others => '0');
signal s845 : std_logic_vector(33 downto 0) := (others => '0');
signal s846 : std_logic_vector(33 downto 0) := (others => '0');
signal s847 : std_logic_vector(33 downto 0) := (others => '0');
signal s848 : std_logic_vector(33 downto 0) := (others => '0');
signal s849 : std_logic_vector(33 downto 0) := (others => '0');
signal s850 : std_logic_vector(33 downto 0) := (others => '0');
signal s851 : std_logic_vector(33 downto 0) := (others => '0');
signal s852 : std_logic_vector(33 downto 0) := (others => '0');
signal s853 : std_logic_vector(33 downto 0) := (others => '0');
signal s854 : std_logic_vector(33 downto 0) := (others => '0');
signal s855 : std_logic_vector(33 downto 0) := (others => '0');
signal s856 : std_logic_vector(33 downto 0) := (others => '0');
signal s857 : std_logic_vector(33 downto 0) := (others => '0');
signal s858 : std_logic_vector(33 downto 0) := (others => '0');
signal s859 : std_logic_vector(33 downto 0) := (others => '0');
signal s860 : std_logic_vector(33 downto 0) := (others => '0');
signal s861 : std_logic_vector(33 downto 0) := (others => '0');
signal s862 : std_logic_vector(33 downto 0) := (others => '0');
signal s863 : std_logic_vector(33 downto 0) := (others => '0');
signal s864 : std_logic_vector(33 downto 0) := (others => '0');
signal s865 : std_logic_vector(33 downto 0) := (others => '0');
signal s866 : std_logic_vector(33 downto 0) := (others => '0');
signal s867 : std_logic_vector(33 downto 0) := (others => '0');
signal s868 : std_logic_vector(33 downto 0) := (others => '0');
signal s869 : std_logic_vector(33 downto 0) := (others => '0');
signal s870 : std_logic_vector(33 downto 0) := (others => '0');
signal s871 : std_logic_vector(33 downto 0) := (others => '0');
signal s872 : std_logic_vector(33 downto 0) := (others => '0');
signal s873 : std_logic_vector(33 downto 0) := (others => '0');
signal s874 : std_logic_vector(33 downto 0) := (others => '0');
signal s875 : std_logic_vector(33 downto 0) := (others => '0');
signal s876 : std_logic_vector(33 downto 0) := (others => '0');
signal s877 : std_logic_vector(33 downto 0) := (others => '0');
signal s878 : std_logic_vector(33 downto 0) := (others => '0');
signal s879 : std_logic_vector(33 downto 0) := (others => '0');
signal s880 : std_logic_vector(33 downto 0) := (others => '0');
signal s881 : std_logic_vector(33 downto 0) := (others => '0');
signal s882 : std_logic_vector(33 downto 0) := (others => '0');
signal s883 : std_logic_vector(33 downto 0) := (others => '0');
signal s884 : std_logic_vector(33 downto 0) := (others => '0');
signal s885 : std_logic_vector(33 downto 0) := (others => '0');
signal s886 : std_logic_vector(33 downto 0) := (others => '0');
signal s887 : std_logic_vector(33 downto 0) := (others => '0');
signal s888 : std_logic_vector(33 downto 0) := (others => '0');
signal s889 : std_logic_vector(33 downto 0) := (others => '0');
signal s890 : std_logic_vector(33 downto 0) := (others => '0');
signal s891 : std_logic_vector(33 downto 0) := (others => '0');
signal s892 : std_logic_vector(33 downto 0) := (others => '0');
signal s893 : std_logic_vector(33 downto 0) := (others => '0');
signal s894 : std_logic_vector(33 downto 0) := (others => '0');
signal s895 : std_logic_vector(33 downto 0) := (others => '0');
signal s896 : std_logic_vector(33 downto 0) := (others => '0');
signal s897 : std_logic_vector(33 downto 0) := (others => '0');
signal s898 : std_logic_vector(33 downto 0) := (others => '0');
signal s899 : std_logic_vector(33 downto 0) := (others => '0');
signal s900 : std_logic_vector(33 downto 0) := (others => '0');
signal s901 : std_logic_vector(33 downto 0) := (others => '0');
signal s902 : std_logic_vector(33 downto 0) := (others => '0');
signal s903 : std_logic_vector(33 downto 0) := (others => '0');
signal s904 : std_logic_vector(33 downto 0) := (others => '0');
signal s905 : std_logic_vector(33 downto 0) := (others => '0');
signal s906 : std_logic_vector(33 downto 0) := (others => '0');
signal s907 : std_logic_vector(33 downto 0) := (others => '0');
signal s908 : std_logic_vector(33 downto 0) := (others => '0');
signal s909 : std_logic_vector(33 downto 0) := (others => '0');
signal s910 : std_logic_vector(33 downto 0) := (others => '0');
signal s911 : std_logic_vector(33 downto 0) := (others => '0');
signal s912 : std_logic_vector(33 downto 0) := (others => '0');
signal s913 : std_logic_vector(33 downto 0) := (others => '0');
signal s914 : std_logic_vector(33 downto 0) := (others => '0');
signal s915 : std_logic_vector(33 downto 0) := (others => '0');
signal s916 : std_logic_vector(33 downto 0) := (others => '0');
signal s917 : std_logic_vector(33 downto 0) := (others => '0');
signal s918 : std_logic_vector(33 downto 0) := (others => '0');
signal s919 : std_logic_vector(33 downto 0) := (others => '0');
signal s920 : std_logic_vector(33 downto 0) := (others => '0');
signal s921 : std_logic_vector(33 downto 0) := (others => '0');
signal s922 : std_logic_vector(33 downto 0) := (others => '0');
signal s923 : std_logic_vector(33 downto 0) := (others => '0');
signal s924 : std_logic_vector(33 downto 0) := (others => '0');
signal s925 : std_logic_vector(33 downto 0) := (others => '0');
signal s926 : std_logic_vector(33 downto 0) := (others => '0');
signal s927 : std_logic_vector(33 downto 0) := (others => '0');
signal s928 : std_logic_vector(33 downto 0) := (others => '0');
signal s929 : std_logic_vector(33 downto 0) := (others => '0');
signal s930 : std_logic_vector(33 downto 0) := (others => '0');
signal s931 : std_logic_vector(33 downto 0) := (others => '0');
signal s932 : std_logic_vector(33 downto 0) := (others => '0');
signal s933 : std_logic_vector(33 downto 0) := (others => '0');
signal s934 : std_logic_vector(33 downto 0) := (others => '0');
signal s935 : std_logic_vector(33 downto 0) := (others => '0');
signal s936 : std_logic_vector(33 downto 0) := (others => '0');
signal s937 : std_logic_vector(33 downto 0) := (others => '0');
signal s938 : std_logic_vector(33 downto 0) := (others => '0');
signal s939 : std_logic_vector(33 downto 0) := (others => '0');
signal s940 : std_logic_vector(33 downto 0) := (others => '0');
signal s941 : std_logic_vector(33 downto 0) := (others => '0');
signal s942 : std_logic_vector(33 downto 0) := (others => '0');
signal s943 : std_logic_vector(33 downto 0) := (others => '0');
signal s944 : std_logic_vector(33 downto 0) := (others => '0');
signal s945 : std_logic_vector(33 downto 0) := (others => '0');
signal s946 : std_logic_vector(33 downto 0) := (others => '0');
signal s947 : std_logic_vector(33 downto 0) := (others => '0');
signal s948 : std_logic_vector(33 downto 0) := (others => '0');
signal s949 : std_logic_vector(33 downto 0) := (others => '0');
signal s950 : std_logic_vector(33 downto 0) := (others => '0');
signal s951 : std_logic_vector(33 downto 0) := (others => '0');
signal s952 : std_logic_vector(33 downto 0) := (others => '0');
signal s953 : std_logic_vector(33 downto 0) := (others => '0');
signal s954 : std_logic_vector(33 downto 0) := (others => '0');
signal s955 : std_logic_vector(33 downto 0) := (others => '0');
signal s956 : std_logic_vector(33 downto 0) := (others => '0');
signal s957 : std_logic_vector(33 downto 0) := (others => '0');
signal s958 : std_logic_vector(33 downto 0) := (others => '0');
signal s959 : std_logic_vector(33 downto 0) := (others => '0');
signal s960 : std_logic_vector(33 downto 0) := (others => '0');
signal s961 : std_logic_vector(33 downto 0) := (others => '0');
signal s962 : std_logic_vector(33 downto 0) := (others => '0');
signal s963 : std_logic_vector(33 downto 0) := (others => '0');
signal s964 : std_logic_vector(33 downto 0) := (others => '0');
signal s965 : std_logic_vector(33 downto 0) := (others => '0');
signal s966 : std_logic_vector(33 downto 0) := (others => '0');
signal s967 : std_logic_vector(33 downto 0) := (others => '0');
signal s968 : std_logic_vector(33 downto 0) := (others => '0');
signal s969 : std_logic_vector(33 downto 0) := (others => '0');
signal s970 : std_logic_vector(33 downto 0) := (others => '0');
signal s971 : std_logic_vector(33 downto 0) := (others => '0');
signal s972 : std_logic_vector(33 downto 0) := (others => '0');
signal s973 : std_logic_vector(33 downto 0) := (others => '0');
signal s974 : std_logic_vector(33 downto 0) := (others => '0');
signal s975 : std_logic_vector(33 downto 0) := (others => '0');
signal s976 : std_logic_vector(33 downto 0) := (others => '0');
signal s977 : std_logic_vector(33 downto 0) := (others => '0');
signal s978 : std_logic_vector(33 downto 0) := (others => '0');
signal s979 : std_logic_vector(33 downto 0) := (others => '0');
signal s980 : std_logic_vector(33 downto 0) := (others => '0');
signal s981 : std_logic_vector(33 downto 0) := (others => '0');
signal s982 : std_logic_vector(33 downto 0) := (others => '0');
signal s983 : std_logic_vector(33 downto 0) := (others => '0');
signal s984 : std_logic_vector(33 downto 0) := (others => '0');
signal s985 : std_logic_vector(33 downto 0) := (others => '0');
signal s986 : std_logic_vector(33 downto 0) := (others => '0');
signal s987 : std_logic_vector(33 downto 0) := (others => '0');
signal s988 : std_logic_vector(33 downto 0) := (others => '0');
signal s989 : std_logic_vector(33 downto 0) := (others => '0');
signal s990 : std_logic_vector(33 downto 0) := (others => '0');
signal s991 : std_logic_vector(33 downto 0) := (others => '0');
signal s992 : std_logic_vector(33 downto 0) := (others => '0');
signal s993 : std_logic_vector(33 downto 0) := (others => '0');
signal s994 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
      s558 <= "0000000000000000000000000000000000";
      s559 <= "0000000000000000000000000000000000";
      s560 <= "0000000000000000000000000000000000";
      s561 <= "0000000000000000000000000000000000";
      s562 <= "0000000000000000000000000000000000";
      s563 <= "0000000000000000000000000000000000";
      s564 <= "0000000000000000000000000000000000";
      s565 <= "0000000000000000000000000000000000";
      s566 <= "0000000000000000000000000000000000";
      s567 <= "0000000000000000000000000000000000";
      s568 <= "0000000000000000000000000000000000";
      s569 <= "0000000000000000000000000000000000";
      s570 <= "0000000000000000000000000000000000";
      s571 <= "0000000000000000000000000000000000";
      s572 <= "0000000000000000000000000000000000";
      s573 <= "0000000000000000000000000000000000";
      s574 <= "0000000000000000000000000000000000";
      s575 <= "0000000000000000000000000000000000";
      s576 <= "0000000000000000000000000000000000";
      s577 <= "0000000000000000000000000000000000";
      s578 <= "0000000000000000000000000000000000";
      s579 <= "0000000000000000000000000000000000";
      s580 <= "0000000000000000000000000000000000";
      s581 <= "0000000000000000000000000000000000";
      s582 <= "0000000000000000000000000000000000";
      s583 <= "0000000000000000000000000000000000";
      s584 <= "0000000000000000000000000000000000";
      s585 <= "0000000000000000000000000000000000";
      s586 <= "0000000000000000000000000000000000";
      s587 <= "0000000000000000000000000000000000";
      s588 <= "0000000000000000000000000000000000";
      s589 <= "0000000000000000000000000000000000";
      s590 <= "0000000000000000000000000000000000";
      s591 <= "0000000000000000000000000000000000";
      s592 <= "0000000000000000000000000000000000";
      s593 <= "0000000000000000000000000000000000";
      s594 <= "0000000000000000000000000000000000";
      s595 <= "0000000000000000000000000000000000";
      s596 <= "0000000000000000000000000000000000";
      s597 <= "0000000000000000000000000000000000";
      s598 <= "0000000000000000000000000000000000";
      s599 <= "0000000000000000000000000000000000";
      s600 <= "0000000000000000000000000000000000";
      s601 <= "0000000000000000000000000000000000";
      s602 <= "0000000000000000000000000000000000";
      s603 <= "0000000000000000000000000000000000";
      s604 <= "0000000000000000000000000000000000";
      s605 <= "0000000000000000000000000000000000";
      s606 <= "0000000000000000000000000000000000";
      s607 <= "0000000000000000000000000000000000";
      s608 <= "0000000000000000000000000000000000";
      s609 <= "0000000000000000000000000000000000";
      s610 <= "0000000000000000000000000000000000";
      s611 <= "0000000000000000000000000000000000";
      s612 <= "0000000000000000000000000000000000";
      s613 <= "0000000000000000000000000000000000";
      s614 <= "0000000000000000000000000000000000";
      s615 <= "0000000000000000000000000000000000";
      s616 <= "0000000000000000000000000000000000";
      s617 <= "0000000000000000000000000000000000";
      s618 <= "0000000000000000000000000000000000";
      s619 <= "0000000000000000000000000000000000";
      s620 <= "0000000000000000000000000000000000";
      s621 <= "0000000000000000000000000000000000";
      s622 <= "0000000000000000000000000000000000";
      s623 <= "0000000000000000000000000000000000";
      s624 <= "0000000000000000000000000000000000";
      s625 <= "0000000000000000000000000000000000";
      s626 <= "0000000000000000000000000000000000";
      s627 <= "0000000000000000000000000000000000";
      s628 <= "0000000000000000000000000000000000";
      s629 <= "0000000000000000000000000000000000";
      s630 <= "0000000000000000000000000000000000";
      s631 <= "0000000000000000000000000000000000";
      s632 <= "0000000000000000000000000000000000";
      s633 <= "0000000000000000000000000000000000";
      s634 <= "0000000000000000000000000000000000";
      s635 <= "0000000000000000000000000000000000";
      s636 <= "0000000000000000000000000000000000";
      s637 <= "0000000000000000000000000000000000";
      s638 <= "0000000000000000000000000000000000";
      s639 <= "0000000000000000000000000000000000";
      s640 <= "0000000000000000000000000000000000";
      s641 <= "0000000000000000000000000000000000";
      s642 <= "0000000000000000000000000000000000";
      s643 <= "0000000000000000000000000000000000";
      s644 <= "0000000000000000000000000000000000";
      s645 <= "0000000000000000000000000000000000";
      s646 <= "0000000000000000000000000000000000";
      s647 <= "0000000000000000000000000000000000";
      s648 <= "0000000000000000000000000000000000";
      s649 <= "0000000000000000000000000000000000";
      s650 <= "0000000000000000000000000000000000";
      s651 <= "0000000000000000000000000000000000";
      s652 <= "0000000000000000000000000000000000";
      s653 <= "0000000000000000000000000000000000";
      s654 <= "0000000000000000000000000000000000";
      s655 <= "0000000000000000000000000000000000";
      s656 <= "0000000000000000000000000000000000";
      s657 <= "0000000000000000000000000000000000";
      s658 <= "0000000000000000000000000000000000";
      s659 <= "0000000000000000000000000000000000";
      s660 <= "0000000000000000000000000000000000";
      s661 <= "0000000000000000000000000000000000";
      s662 <= "0000000000000000000000000000000000";
      s663 <= "0000000000000000000000000000000000";
      s664 <= "0000000000000000000000000000000000";
      s665 <= "0000000000000000000000000000000000";
      s666 <= "0000000000000000000000000000000000";
      s667 <= "0000000000000000000000000000000000";
      s668 <= "0000000000000000000000000000000000";
      s669 <= "0000000000000000000000000000000000";
      s670 <= "0000000000000000000000000000000000";
      s671 <= "0000000000000000000000000000000000";
      s672 <= "0000000000000000000000000000000000";
      s673 <= "0000000000000000000000000000000000";
      s674 <= "0000000000000000000000000000000000";
      s675 <= "0000000000000000000000000000000000";
      s676 <= "0000000000000000000000000000000000";
      s677 <= "0000000000000000000000000000000000";
      s678 <= "0000000000000000000000000000000000";
      s679 <= "0000000000000000000000000000000000";
      s680 <= "0000000000000000000000000000000000";
      s681 <= "0000000000000000000000000000000000";
      s682 <= "0000000000000000000000000000000000";
      s683 <= "0000000000000000000000000000000000";
      s684 <= "0000000000000000000000000000000000";
      s685 <= "0000000000000000000000000000000000";
      s686 <= "0000000000000000000000000000000000";
      s687 <= "0000000000000000000000000000000000";
      s688 <= "0000000000000000000000000000000000";
      s689 <= "0000000000000000000000000000000000";
      s690 <= "0000000000000000000000000000000000";
      s691 <= "0000000000000000000000000000000000";
      s692 <= "0000000000000000000000000000000000";
      s693 <= "0000000000000000000000000000000000";
      s694 <= "0000000000000000000000000000000000";
      s695 <= "0000000000000000000000000000000000";
      s696 <= "0000000000000000000000000000000000";
      s697 <= "0000000000000000000000000000000000";
      s698 <= "0000000000000000000000000000000000";
      s699 <= "0000000000000000000000000000000000";
      s700 <= "0000000000000000000000000000000000";
      s701 <= "0000000000000000000000000000000000";
      s702 <= "0000000000000000000000000000000000";
      s703 <= "0000000000000000000000000000000000";
      s704 <= "0000000000000000000000000000000000";
      s705 <= "0000000000000000000000000000000000";
      s706 <= "0000000000000000000000000000000000";
      s707 <= "0000000000000000000000000000000000";
      s708 <= "0000000000000000000000000000000000";
      s709 <= "0000000000000000000000000000000000";
      s710 <= "0000000000000000000000000000000000";
      s711 <= "0000000000000000000000000000000000";
      s712 <= "0000000000000000000000000000000000";
      s713 <= "0000000000000000000000000000000000";
      s714 <= "0000000000000000000000000000000000";
      s715 <= "0000000000000000000000000000000000";
      s716 <= "0000000000000000000000000000000000";
      s717 <= "0000000000000000000000000000000000";
      s718 <= "0000000000000000000000000000000000";
      s719 <= "0000000000000000000000000000000000";
      s720 <= "0000000000000000000000000000000000";
      s721 <= "0000000000000000000000000000000000";
      s722 <= "0000000000000000000000000000000000";
      s723 <= "0000000000000000000000000000000000";
      s724 <= "0000000000000000000000000000000000";
      s725 <= "0000000000000000000000000000000000";
      s726 <= "0000000000000000000000000000000000";
      s727 <= "0000000000000000000000000000000000";
      s728 <= "0000000000000000000000000000000000";
      s729 <= "0000000000000000000000000000000000";
      s730 <= "0000000000000000000000000000000000";
      s731 <= "0000000000000000000000000000000000";
      s732 <= "0000000000000000000000000000000000";
      s733 <= "0000000000000000000000000000000000";
      s734 <= "0000000000000000000000000000000000";
      s735 <= "0000000000000000000000000000000000";
      s736 <= "0000000000000000000000000000000000";
      s737 <= "0000000000000000000000000000000000";
      s738 <= "0000000000000000000000000000000000";
      s739 <= "0000000000000000000000000000000000";
      s740 <= "0000000000000000000000000000000000";
      s741 <= "0000000000000000000000000000000000";
      s742 <= "0000000000000000000000000000000000";
      s743 <= "0000000000000000000000000000000000";
      s744 <= "0000000000000000000000000000000000";
      s745 <= "0000000000000000000000000000000000";
      s746 <= "0000000000000000000000000000000000";
      s747 <= "0000000000000000000000000000000000";
      s748 <= "0000000000000000000000000000000000";
      s749 <= "0000000000000000000000000000000000";
      s750 <= "0000000000000000000000000000000000";
      s751 <= "0000000000000000000000000000000000";
      s752 <= "0000000000000000000000000000000000";
      s753 <= "0000000000000000000000000000000000";
      s754 <= "0000000000000000000000000000000000";
      s755 <= "0000000000000000000000000000000000";
      s756 <= "0000000000000000000000000000000000";
      s757 <= "0000000000000000000000000000000000";
      s758 <= "0000000000000000000000000000000000";
      s759 <= "0000000000000000000000000000000000";
      s760 <= "0000000000000000000000000000000000";
      s761 <= "0000000000000000000000000000000000";
      s762 <= "0000000000000000000000000000000000";
      s763 <= "0000000000000000000000000000000000";
      s764 <= "0000000000000000000000000000000000";
      s765 <= "0000000000000000000000000000000000";
      s766 <= "0000000000000000000000000000000000";
      s767 <= "0000000000000000000000000000000000";
      s768 <= "0000000000000000000000000000000000";
      s769 <= "0000000000000000000000000000000000";
      s770 <= "0000000000000000000000000000000000";
      s771 <= "0000000000000000000000000000000000";
      s772 <= "0000000000000000000000000000000000";
      s773 <= "0000000000000000000000000000000000";
      s774 <= "0000000000000000000000000000000000";
      s775 <= "0000000000000000000000000000000000";
      s776 <= "0000000000000000000000000000000000";
      s777 <= "0000000000000000000000000000000000";
      s778 <= "0000000000000000000000000000000000";
      s779 <= "0000000000000000000000000000000000";
      s780 <= "0000000000000000000000000000000000";
      s781 <= "0000000000000000000000000000000000";
      s782 <= "0000000000000000000000000000000000";
      s783 <= "0000000000000000000000000000000000";
      s784 <= "0000000000000000000000000000000000";
      s785 <= "0000000000000000000000000000000000";
      s786 <= "0000000000000000000000000000000000";
      s787 <= "0000000000000000000000000000000000";
      s788 <= "0000000000000000000000000000000000";
      s789 <= "0000000000000000000000000000000000";
      s790 <= "0000000000000000000000000000000000";
      s791 <= "0000000000000000000000000000000000";
      s792 <= "0000000000000000000000000000000000";
      s793 <= "0000000000000000000000000000000000";
      s794 <= "0000000000000000000000000000000000";
      s795 <= "0000000000000000000000000000000000";
      s796 <= "0000000000000000000000000000000000";
      s797 <= "0000000000000000000000000000000000";
      s798 <= "0000000000000000000000000000000000";
      s799 <= "0000000000000000000000000000000000";
      s800 <= "0000000000000000000000000000000000";
      s801 <= "0000000000000000000000000000000000";
      s802 <= "0000000000000000000000000000000000";
      s803 <= "0000000000000000000000000000000000";
      s804 <= "0000000000000000000000000000000000";
      s805 <= "0000000000000000000000000000000000";
      s806 <= "0000000000000000000000000000000000";
      s807 <= "0000000000000000000000000000000000";
      s808 <= "0000000000000000000000000000000000";
      s809 <= "0000000000000000000000000000000000";
      s810 <= "0000000000000000000000000000000000";
      s811 <= "0000000000000000000000000000000000";
      s812 <= "0000000000000000000000000000000000";
      s813 <= "0000000000000000000000000000000000";
      s814 <= "0000000000000000000000000000000000";
      s815 <= "0000000000000000000000000000000000";
      s816 <= "0000000000000000000000000000000000";
      s817 <= "0000000000000000000000000000000000";
      s818 <= "0000000000000000000000000000000000";
      s819 <= "0000000000000000000000000000000000";
      s820 <= "0000000000000000000000000000000000";
      s821 <= "0000000000000000000000000000000000";
      s822 <= "0000000000000000000000000000000000";
      s823 <= "0000000000000000000000000000000000";
      s824 <= "0000000000000000000000000000000000";
      s825 <= "0000000000000000000000000000000000";
      s826 <= "0000000000000000000000000000000000";
      s827 <= "0000000000000000000000000000000000";
      s828 <= "0000000000000000000000000000000000";
      s829 <= "0000000000000000000000000000000000";
      s830 <= "0000000000000000000000000000000000";
      s831 <= "0000000000000000000000000000000000";
      s832 <= "0000000000000000000000000000000000";
      s833 <= "0000000000000000000000000000000000";
      s834 <= "0000000000000000000000000000000000";
      s835 <= "0000000000000000000000000000000000";
      s836 <= "0000000000000000000000000000000000";
      s837 <= "0000000000000000000000000000000000";
      s838 <= "0000000000000000000000000000000000";
      s839 <= "0000000000000000000000000000000000";
      s840 <= "0000000000000000000000000000000000";
      s841 <= "0000000000000000000000000000000000";
      s842 <= "0000000000000000000000000000000000";
      s843 <= "0000000000000000000000000000000000";
      s844 <= "0000000000000000000000000000000000";
      s845 <= "0000000000000000000000000000000000";
      s846 <= "0000000000000000000000000000000000";
      s847 <= "0000000000000000000000000000000000";
      s848 <= "0000000000000000000000000000000000";
      s849 <= "0000000000000000000000000000000000";
      s850 <= "0000000000000000000000000000000000";
      s851 <= "0000000000000000000000000000000000";
      s852 <= "0000000000000000000000000000000000";
      s853 <= "0000000000000000000000000000000000";
      s854 <= "0000000000000000000000000000000000";
      s855 <= "0000000000000000000000000000000000";
      s856 <= "0000000000000000000000000000000000";
      s857 <= "0000000000000000000000000000000000";
      s858 <= "0000000000000000000000000000000000";
      s859 <= "0000000000000000000000000000000000";
      s860 <= "0000000000000000000000000000000000";
      s861 <= "0000000000000000000000000000000000";
      s862 <= "0000000000000000000000000000000000";
      s863 <= "0000000000000000000000000000000000";
      s864 <= "0000000000000000000000000000000000";
      s865 <= "0000000000000000000000000000000000";
      s866 <= "0000000000000000000000000000000000";
      s867 <= "0000000000000000000000000000000000";
      s868 <= "0000000000000000000000000000000000";
      s869 <= "0000000000000000000000000000000000";
      s870 <= "0000000000000000000000000000000000";
      s871 <= "0000000000000000000000000000000000";
      s872 <= "0000000000000000000000000000000000";
      s873 <= "0000000000000000000000000000000000";
      s874 <= "0000000000000000000000000000000000";
      s875 <= "0000000000000000000000000000000000";
      s876 <= "0000000000000000000000000000000000";
      s877 <= "0000000000000000000000000000000000";
      s878 <= "0000000000000000000000000000000000";
      s879 <= "0000000000000000000000000000000000";
      s880 <= "0000000000000000000000000000000000";
      s881 <= "0000000000000000000000000000000000";
      s882 <= "0000000000000000000000000000000000";
      s883 <= "0000000000000000000000000000000000";
      s884 <= "0000000000000000000000000000000000";
      s885 <= "0000000000000000000000000000000000";
      s886 <= "0000000000000000000000000000000000";
      s887 <= "0000000000000000000000000000000000";
      s888 <= "0000000000000000000000000000000000";
      s889 <= "0000000000000000000000000000000000";
      s890 <= "0000000000000000000000000000000000";
      s891 <= "0000000000000000000000000000000000";
      s892 <= "0000000000000000000000000000000000";
      s893 <= "0000000000000000000000000000000000";
      s894 <= "0000000000000000000000000000000000";
      s895 <= "0000000000000000000000000000000000";
      s896 <= "0000000000000000000000000000000000";
      s897 <= "0000000000000000000000000000000000";
      s898 <= "0000000000000000000000000000000000";
      s899 <= "0000000000000000000000000000000000";
      s900 <= "0000000000000000000000000000000000";
      s901 <= "0000000000000000000000000000000000";
      s902 <= "0000000000000000000000000000000000";
      s903 <= "0000000000000000000000000000000000";
      s904 <= "0000000000000000000000000000000000";
      s905 <= "0000000000000000000000000000000000";
      s906 <= "0000000000000000000000000000000000";
      s907 <= "0000000000000000000000000000000000";
      s908 <= "0000000000000000000000000000000000";
      s909 <= "0000000000000000000000000000000000";
      s910 <= "0000000000000000000000000000000000";
      s911 <= "0000000000000000000000000000000000";
      s912 <= "0000000000000000000000000000000000";
      s913 <= "0000000000000000000000000000000000";
      s914 <= "0000000000000000000000000000000000";
      s915 <= "0000000000000000000000000000000000";
      s916 <= "0000000000000000000000000000000000";
      s917 <= "0000000000000000000000000000000000";
      s918 <= "0000000000000000000000000000000000";
      s919 <= "0000000000000000000000000000000000";
      s920 <= "0000000000000000000000000000000000";
      s921 <= "0000000000000000000000000000000000";
      s922 <= "0000000000000000000000000000000000";
      s923 <= "0000000000000000000000000000000000";
      s924 <= "0000000000000000000000000000000000";
      s925 <= "0000000000000000000000000000000000";
      s926 <= "0000000000000000000000000000000000";
      s927 <= "0000000000000000000000000000000000";
      s928 <= "0000000000000000000000000000000000";
      s929 <= "0000000000000000000000000000000000";
      s930 <= "0000000000000000000000000000000000";
      s931 <= "0000000000000000000000000000000000";
      s932 <= "0000000000000000000000000000000000";
      s933 <= "0000000000000000000000000000000000";
      s934 <= "0000000000000000000000000000000000";
      s935 <= "0000000000000000000000000000000000";
      s936 <= "0000000000000000000000000000000000";
      s937 <= "0000000000000000000000000000000000";
      s938 <= "0000000000000000000000000000000000";
      s939 <= "0000000000000000000000000000000000";
      s940 <= "0000000000000000000000000000000000";
      s941 <= "0000000000000000000000000000000000";
      s942 <= "0000000000000000000000000000000000";
      s943 <= "0000000000000000000000000000000000";
      s944 <= "0000000000000000000000000000000000";
      s945 <= "0000000000000000000000000000000000";
      s946 <= "0000000000000000000000000000000000";
      s947 <= "0000000000000000000000000000000000";
      s948 <= "0000000000000000000000000000000000";
      s949 <= "0000000000000000000000000000000000";
      s950 <= "0000000000000000000000000000000000";
      s951 <= "0000000000000000000000000000000000";
      s952 <= "0000000000000000000000000000000000";
      s953 <= "0000000000000000000000000000000000";
      s954 <= "0000000000000000000000000000000000";
      s955 <= "0000000000000000000000000000000000";
      s956 <= "0000000000000000000000000000000000";
      s957 <= "0000000000000000000000000000000000";
      s958 <= "0000000000000000000000000000000000";
      s959 <= "0000000000000000000000000000000000";
      s960 <= "0000000000000000000000000000000000";
      s961 <= "0000000000000000000000000000000000";
      s962 <= "0000000000000000000000000000000000";
      s963 <= "0000000000000000000000000000000000";
      s964 <= "0000000000000000000000000000000000";
      s965 <= "0000000000000000000000000000000000";
      s966 <= "0000000000000000000000000000000000";
      s967 <= "0000000000000000000000000000000000";
      s968 <= "0000000000000000000000000000000000";
      s969 <= "0000000000000000000000000000000000";
      s970 <= "0000000000000000000000000000000000";
      s971 <= "0000000000000000000000000000000000";
      s972 <= "0000000000000000000000000000000000";
      s973 <= "0000000000000000000000000000000000";
      s974 <= "0000000000000000000000000000000000";
      s975 <= "0000000000000000000000000000000000";
      s976 <= "0000000000000000000000000000000000";
      s977 <= "0000000000000000000000000000000000";
      s978 <= "0000000000000000000000000000000000";
      s979 <= "0000000000000000000000000000000000";
      s980 <= "0000000000000000000000000000000000";
      s981 <= "0000000000000000000000000000000000";
      s982 <= "0000000000000000000000000000000000";
      s983 <= "0000000000000000000000000000000000";
      s984 <= "0000000000000000000000000000000000";
      s985 <= "0000000000000000000000000000000000";
      s986 <= "0000000000000000000000000000000000";
      s987 <= "0000000000000000000000000000000000";
      s988 <= "0000000000000000000000000000000000";
      s989 <= "0000000000000000000000000000000000";
      s990 <= "0000000000000000000000000000000000";
      s991 <= "0000000000000000000000000000000000";
      s992 <= "0000000000000000000000000000000000";
      s993 <= "0000000000000000000000000000000000";
      s994 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      s558 <= s557;
      s559 <= s558;
      s560 <= s559;
      s561 <= s560;
      s562 <= s561;
      s563 <= s562;
      s564 <= s563;
      s565 <= s564;
      s566 <= s565;
      s567 <= s566;
      s568 <= s567;
      s569 <= s568;
      s570 <= s569;
      s571 <= s570;
      s572 <= s571;
      s573 <= s572;
      s574 <= s573;
      s575 <= s574;
      s576 <= s575;
      s577 <= s576;
      s578 <= s577;
      s579 <= s578;
      s580 <= s579;
      s581 <= s580;
      s582 <= s581;
      s583 <= s582;
      s584 <= s583;
      s585 <= s584;
      s586 <= s585;
      s587 <= s586;
      s588 <= s587;
      s589 <= s588;
      s590 <= s589;
      s591 <= s590;
      s592 <= s591;
      s593 <= s592;
      s594 <= s593;
      s595 <= s594;
      s596 <= s595;
      s597 <= s596;
      s598 <= s597;
      s599 <= s598;
      s600 <= s599;
      s601 <= s600;
      s602 <= s601;
      s603 <= s602;
      s604 <= s603;
      s605 <= s604;
      s606 <= s605;
      s607 <= s606;
      s608 <= s607;
      s609 <= s608;
      s610 <= s609;
      s611 <= s610;
      s612 <= s611;
      s613 <= s612;
      s614 <= s613;
      s615 <= s614;
      s616 <= s615;
      s617 <= s616;
      s618 <= s617;
      s619 <= s618;
      s620 <= s619;
      s621 <= s620;
      s622 <= s621;
      s623 <= s622;
      s624 <= s623;
      s625 <= s624;
      s626 <= s625;
      s627 <= s626;
      s628 <= s627;
      s629 <= s628;
      s630 <= s629;
      s631 <= s630;
      s632 <= s631;
      s633 <= s632;
      s634 <= s633;
      s635 <= s634;
      s636 <= s635;
      s637 <= s636;
      s638 <= s637;
      s639 <= s638;
      s640 <= s639;
      s641 <= s640;
      s642 <= s641;
      s643 <= s642;
      s644 <= s643;
      s645 <= s644;
      s646 <= s645;
      s647 <= s646;
      s648 <= s647;
      s649 <= s648;
      s650 <= s649;
      s651 <= s650;
      s652 <= s651;
      s653 <= s652;
      s654 <= s653;
      s655 <= s654;
      s656 <= s655;
      s657 <= s656;
      s658 <= s657;
      s659 <= s658;
      s660 <= s659;
      s661 <= s660;
      s662 <= s661;
      s663 <= s662;
      s664 <= s663;
      s665 <= s664;
      s666 <= s665;
      s667 <= s666;
      s668 <= s667;
      s669 <= s668;
      s670 <= s669;
      s671 <= s670;
      s672 <= s671;
      s673 <= s672;
      s674 <= s673;
      s675 <= s674;
      s676 <= s675;
      s677 <= s676;
      s678 <= s677;
      s679 <= s678;
      s680 <= s679;
      s681 <= s680;
      s682 <= s681;
      s683 <= s682;
      s684 <= s683;
      s685 <= s684;
      s686 <= s685;
      s687 <= s686;
      s688 <= s687;
      s689 <= s688;
      s690 <= s689;
      s691 <= s690;
      s692 <= s691;
      s693 <= s692;
      s694 <= s693;
      s695 <= s694;
      s696 <= s695;
      s697 <= s696;
      s698 <= s697;
      s699 <= s698;
      s700 <= s699;
      s701 <= s700;
      s702 <= s701;
      s703 <= s702;
      s704 <= s703;
      s705 <= s704;
      s706 <= s705;
      s707 <= s706;
      s708 <= s707;
      s709 <= s708;
      s710 <= s709;
      s711 <= s710;
      s712 <= s711;
      s713 <= s712;
      s714 <= s713;
      s715 <= s714;
      s716 <= s715;
      s717 <= s716;
      s718 <= s717;
      s719 <= s718;
      s720 <= s719;
      s721 <= s720;
      s722 <= s721;
      s723 <= s722;
      s724 <= s723;
      s725 <= s724;
      s726 <= s725;
      s727 <= s726;
      s728 <= s727;
      s729 <= s728;
      s730 <= s729;
      s731 <= s730;
      s732 <= s731;
      s733 <= s732;
      s734 <= s733;
      s735 <= s734;
      s736 <= s735;
      s737 <= s736;
      s738 <= s737;
      s739 <= s738;
      s740 <= s739;
      s741 <= s740;
      s742 <= s741;
      s743 <= s742;
      s744 <= s743;
      s745 <= s744;
      s746 <= s745;
      s747 <= s746;
      s748 <= s747;
      s749 <= s748;
      s750 <= s749;
      s751 <= s750;
      s752 <= s751;
      s753 <= s752;
      s754 <= s753;
      s755 <= s754;
      s756 <= s755;
      s757 <= s756;
      s758 <= s757;
      s759 <= s758;
      s760 <= s759;
      s761 <= s760;
      s762 <= s761;
      s763 <= s762;
      s764 <= s763;
      s765 <= s764;
      s766 <= s765;
      s767 <= s766;
      s768 <= s767;
      s769 <= s768;
      s770 <= s769;
      s771 <= s770;
      s772 <= s771;
      s773 <= s772;
      s774 <= s773;
      s775 <= s774;
      s776 <= s775;
      s777 <= s776;
      s778 <= s777;
      s779 <= s778;
      s780 <= s779;
      s781 <= s780;
      s782 <= s781;
      s783 <= s782;
      s784 <= s783;
      s785 <= s784;
      s786 <= s785;
      s787 <= s786;
      s788 <= s787;
      s789 <= s788;
      s790 <= s789;
      s791 <= s790;
      s792 <= s791;
      s793 <= s792;
      s794 <= s793;
      s795 <= s794;
      s796 <= s795;
      s797 <= s796;
      s798 <= s797;
      s799 <= s798;
      s800 <= s799;
      s801 <= s800;
      s802 <= s801;
      s803 <= s802;
      s804 <= s803;
      s805 <= s804;
      s806 <= s805;
      s807 <= s806;
      s808 <= s807;
      s809 <= s808;
      s810 <= s809;
      s811 <= s810;
      s812 <= s811;
      s813 <= s812;
      s814 <= s813;
      s815 <= s814;
      s816 <= s815;
      s817 <= s816;
      s818 <= s817;
      s819 <= s818;
      s820 <= s819;
      s821 <= s820;
      s822 <= s821;
      s823 <= s822;
      s824 <= s823;
      s825 <= s824;
      s826 <= s825;
      s827 <= s826;
      s828 <= s827;
      s829 <= s828;
      s830 <= s829;
      s831 <= s830;
      s832 <= s831;
      s833 <= s832;
      s834 <= s833;
      s835 <= s834;
      s836 <= s835;
      s837 <= s836;
      s838 <= s837;
      s839 <= s838;
      s840 <= s839;
      s841 <= s840;
      s842 <= s841;
      s843 <= s842;
      s844 <= s843;
      s845 <= s844;
      s846 <= s845;
      s847 <= s846;
      s848 <= s847;
      s849 <= s848;
      s850 <= s849;
      s851 <= s850;
      s852 <= s851;
      s853 <= s852;
      s854 <= s853;
      s855 <= s854;
      s856 <= s855;
      s857 <= s856;
      s858 <= s857;
      s859 <= s858;
      s860 <= s859;
      s861 <= s860;
      s862 <= s861;
      s863 <= s862;
      s864 <= s863;
      s865 <= s864;
      s866 <= s865;
      s867 <= s866;
      s868 <= s867;
      s869 <= s868;
      s870 <= s869;
      s871 <= s870;
      s872 <= s871;
      s873 <= s872;
      s874 <= s873;
      s875 <= s874;
      s876 <= s875;
      s877 <= s876;
      s878 <= s877;
      s879 <= s878;
      s880 <= s879;
      s881 <= s880;
      s882 <= s881;
      s883 <= s882;
      s884 <= s883;
      s885 <= s884;
      s886 <= s885;
      s887 <= s886;
      s888 <= s887;
      s889 <= s888;
      s890 <= s889;
      s891 <= s890;
      s892 <= s891;
      s893 <= s892;
      s894 <= s893;
      s895 <= s894;
      s896 <= s895;
      s897 <= s896;
      s898 <= s897;
      s899 <= s898;
      s900 <= s899;
      s901 <= s900;
      s902 <= s901;
      s903 <= s902;
      s904 <= s903;
      s905 <= s904;
      s906 <= s905;
      s907 <= s906;
      s908 <= s907;
      s909 <= s908;
      s910 <= s909;
      s911 <= s910;
      s912 <= s911;
      s913 <= s912;
      s914 <= s913;
      s915 <= s914;
      s916 <= s915;
      s917 <= s916;
      s918 <= s917;
      s919 <= s918;
      s920 <= s919;
      s921 <= s920;
      s922 <= s921;
      s923 <= s922;
      s924 <= s923;
      s925 <= s924;
      s926 <= s925;
      s927 <= s926;
      s928 <= s927;
      s929 <= s928;
      s930 <= s929;
      s931 <= s930;
      s932 <= s931;
      s933 <= s932;
      s934 <= s933;
      s935 <= s934;
      s936 <= s935;
      s937 <= s936;
      s938 <= s937;
      s939 <= s938;
      s940 <= s939;
      s941 <= s940;
      s942 <= s941;
      s943 <= s942;
      s944 <= s943;
      s945 <= s944;
      s946 <= s945;
      s947 <= s946;
      s948 <= s947;
      s949 <= s948;
      s950 <= s949;
      s951 <= s950;
      s952 <= s951;
      s953 <= s952;
      s954 <= s953;
      s955 <= s954;
      s956 <= s955;
      s957 <= s956;
      s958 <= s957;
      s959 <= s958;
      s960 <= s959;
      s961 <= s960;
      s962 <= s961;
      s963 <= s962;
      s964 <= s963;
      s965 <= s964;
      s966 <= s965;
      s967 <= s966;
      s968 <= s967;
      s969 <= s968;
      s970 <= s969;
      s971 <= s970;
      s972 <= s971;
      s973 <= s972;
      s974 <= s973;
      s975 <= s974;
      s976 <= s975;
      s977 <= s976;
      s978 <= s977;
      s979 <= s978;
      s980 <= s979;
      s981 <= s980;
      s982 <= s981;
      s983 <= s982;
      s984 <= s983;
      s985 <= s984;
      s986 <= s985;
      s987 <= s986;
      s988 <= s987;
      s989 <= s988;
      s990 <= s989;
      s991 <= s990;
      s992 <= s991;
      s993 <= s992;
      s994 <= s993;
      Y <= s994;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1056_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1056 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1056_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1056_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
signal s558 : std_logic_vector(33 downto 0) := (others => '0');
signal s559 : std_logic_vector(33 downto 0) := (others => '0');
signal s560 : std_logic_vector(33 downto 0) := (others => '0');
signal s561 : std_logic_vector(33 downto 0) := (others => '0');
signal s562 : std_logic_vector(33 downto 0) := (others => '0');
signal s563 : std_logic_vector(33 downto 0) := (others => '0');
signal s564 : std_logic_vector(33 downto 0) := (others => '0');
signal s565 : std_logic_vector(33 downto 0) := (others => '0');
signal s566 : std_logic_vector(33 downto 0) := (others => '0');
signal s567 : std_logic_vector(33 downto 0) := (others => '0');
signal s568 : std_logic_vector(33 downto 0) := (others => '0');
signal s569 : std_logic_vector(33 downto 0) := (others => '0');
signal s570 : std_logic_vector(33 downto 0) := (others => '0');
signal s571 : std_logic_vector(33 downto 0) := (others => '0');
signal s572 : std_logic_vector(33 downto 0) := (others => '0');
signal s573 : std_logic_vector(33 downto 0) := (others => '0');
signal s574 : std_logic_vector(33 downto 0) := (others => '0');
signal s575 : std_logic_vector(33 downto 0) := (others => '0');
signal s576 : std_logic_vector(33 downto 0) := (others => '0');
signal s577 : std_logic_vector(33 downto 0) := (others => '0');
signal s578 : std_logic_vector(33 downto 0) := (others => '0');
signal s579 : std_logic_vector(33 downto 0) := (others => '0');
signal s580 : std_logic_vector(33 downto 0) := (others => '0');
signal s581 : std_logic_vector(33 downto 0) := (others => '0');
signal s582 : std_logic_vector(33 downto 0) := (others => '0');
signal s583 : std_logic_vector(33 downto 0) := (others => '0');
signal s584 : std_logic_vector(33 downto 0) := (others => '0');
signal s585 : std_logic_vector(33 downto 0) := (others => '0');
signal s586 : std_logic_vector(33 downto 0) := (others => '0');
signal s587 : std_logic_vector(33 downto 0) := (others => '0');
signal s588 : std_logic_vector(33 downto 0) := (others => '0');
signal s589 : std_logic_vector(33 downto 0) := (others => '0');
signal s590 : std_logic_vector(33 downto 0) := (others => '0');
signal s591 : std_logic_vector(33 downto 0) := (others => '0');
signal s592 : std_logic_vector(33 downto 0) := (others => '0');
signal s593 : std_logic_vector(33 downto 0) := (others => '0');
signal s594 : std_logic_vector(33 downto 0) := (others => '0');
signal s595 : std_logic_vector(33 downto 0) := (others => '0');
signal s596 : std_logic_vector(33 downto 0) := (others => '0');
signal s597 : std_logic_vector(33 downto 0) := (others => '0');
signal s598 : std_logic_vector(33 downto 0) := (others => '0');
signal s599 : std_logic_vector(33 downto 0) := (others => '0');
signal s600 : std_logic_vector(33 downto 0) := (others => '0');
signal s601 : std_logic_vector(33 downto 0) := (others => '0');
signal s602 : std_logic_vector(33 downto 0) := (others => '0');
signal s603 : std_logic_vector(33 downto 0) := (others => '0');
signal s604 : std_logic_vector(33 downto 0) := (others => '0');
signal s605 : std_logic_vector(33 downto 0) := (others => '0');
signal s606 : std_logic_vector(33 downto 0) := (others => '0');
signal s607 : std_logic_vector(33 downto 0) := (others => '0');
signal s608 : std_logic_vector(33 downto 0) := (others => '0');
signal s609 : std_logic_vector(33 downto 0) := (others => '0');
signal s610 : std_logic_vector(33 downto 0) := (others => '0');
signal s611 : std_logic_vector(33 downto 0) := (others => '0');
signal s612 : std_logic_vector(33 downto 0) := (others => '0');
signal s613 : std_logic_vector(33 downto 0) := (others => '0');
signal s614 : std_logic_vector(33 downto 0) := (others => '0');
signal s615 : std_logic_vector(33 downto 0) := (others => '0');
signal s616 : std_logic_vector(33 downto 0) := (others => '0');
signal s617 : std_logic_vector(33 downto 0) := (others => '0');
signal s618 : std_logic_vector(33 downto 0) := (others => '0');
signal s619 : std_logic_vector(33 downto 0) := (others => '0');
signal s620 : std_logic_vector(33 downto 0) := (others => '0');
signal s621 : std_logic_vector(33 downto 0) := (others => '0');
signal s622 : std_logic_vector(33 downto 0) := (others => '0');
signal s623 : std_logic_vector(33 downto 0) := (others => '0');
signal s624 : std_logic_vector(33 downto 0) := (others => '0');
signal s625 : std_logic_vector(33 downto 0) := (others => '0');
signal s626 : std_logic_vector(33 downto 0) := (others => '0');
signal s627 : std_logic_vector(33 downto 0) := (others => '0');
signal s628 : std_logic_vector(33 downto 0) := (others => '0');
signal s629 : std_logic_vector(33 downto 0) := (others => '0');
signal s630 : std_logic_vector(33 downto 0) := (others => '0');
signal s631 : std_logic_vector(33 downto 0) := (others => '0');
signal s632 : std_logic_vector(33 downto 0) := (others => '0');
signal s633 : std_logic_vector(33 downto 0) := (others => '0');
signal s634 : std_logic_vector(33 downto 0) := (others => '0');
signal s635 : std_logic_vector(33 downto 0) := (others => '0');
signal s636 : std_logic_vector(33 downto 0) := (others => '0');
signal s637 : std_logic_vector(33 downto 0) := (others => '0');
signal s638 : std_logic_vector(33 downto 0) := (others => '0');
signal s639 : std_logic_vector(33 downto 0) := (others => '0');
signal s640 : std_logic_vector(33 downto 0) := (others => '0');
signal s641 : std_logic_vector(33 downto 0) := (others => '0');
signal s642 : std_logic_vector(33 downto 0) := (others => '0');
signal s643 : std_logic_vector(33 downto 0) := (others => '0');
signal s644 : std_logic_vector(33 downto 0) := (others => '0');
signal s645 : std_logic_vector(33 downto 0) := (others => '0');
signal s646 : std_logic_vector(33 downto 0) := (others => '0');
signal s647 : std_logic_vector(33 downto 0) := (others => '0');
signal s648 : std_logic_vector(33 downto 0) := (others => '0');
signal s649 : std_logic_vector(33 downto 0) := (others => '0');
signal s650 : std_logic_vector(33 downto 0) := (others => '0');
signal s651 : std_logic_vector(33 downto 0) := (others => '0');
signal s652 : std_logic_vector(33 downto 0) := (others => '0');
signal s653 : std_logic_vector(33 downto 0) := (others => '0');
signal s654 : std_logic_vector(33 downto 0) := (others => '0');
signal s655 : std_logic_vector(33 downto 0) := (others => '0');
signal s656 : std_logic_vector(33 downto 0) := (others => '0');
signal s657 : std_logic_vector(33 downto 0) := (others => '0');
signal s658 : std_logic_vector(33 downto 0) := (others => '0');
signal s659 : std_logic_vector(33 downto 0) := (others => '0');
signal s660 : std_logic_vector(33 downto 0) := (others => '0');
signal s661 : std_logic_vector(33 downto 0) := (others => '0');
signal s662 : std_logic_vector(33 downto 0) := (others => '0');
signal s663 : std_logic_vector(33 downto 0) := (others => '0');
signal s664 : std_logic_vector(33 downto 0) := (others => '0');
signal s665 : std_logic_vector(33 downto 0) := (others => '0');
signal s666 : std_logic_vector(33 downto 0) := (others => '0');
signal s667 : std_logic_vector(33 downto 0) := (others => '0');
signal s668 : std_logic_vector(33 downto 0) := (others => '0');
signal s669 : std_logic_vector(33 downto 0) := (others => '0');
signal s670 : std_logic_vector(33 downto 0) := (others => '0');
signal s671 : std_logic_vector(33 downto 0) := (others => '0');
signal s672 : std_logic_vector(33 downto 0) := (others => '0');
signal s673 : std_logic_vector(33 downto 0) := (others => '0');
signal s674 : std_logic_vector(33 downto 0) := (others => '0');
signal s675 : std_logic_vector(33 downto 0) := (others => '0');
signal s676 : std_logic_vector(33 downto 0) := (others => '0');
signal s677 : std_logic_vector(33 downto 0) := (others => '0');
signal s678 : std_logic_vector(33 downto 0) := (others => '0');
signal s679 : std_logic_vector(33 downto 0) := (others => '0');
signal s680 : std_logic_vector(33 downto 0) := (others => '0');
signal s681 : std_logic_vector(33 downto 0) := (others => '0');
signal s682 : std_logic_vector(33 downto 0) := (others => '0');
signal s683 : std_logic_vector(33 downto 0) := (others => '0');
signal s684 : std_logic_vector(33 downto 0) := (others => '0');
signal s685 : std_logic_vector(33 downto 0) := (others => '0');
signal s686 : std_logic_vector(33 downto 0) := (others => '0');
signal s687 : std_logic_vector(33 downto 0) := (others => '0');
signal s688 : std_logic_vector(33 downto 0) := (others => '0');
signal s689 : std_logic_vector(33 downto 0) := (others => '0');
signal s690 : std_logic_vector(33 downto 0) := (others => '0');
signal s691 : std_logic_vector(33 downto 0) := (others => '0');
signal s692 : std_logic_vector(33 downto 0) := (others => '0');
signal s693 : std_logic_vector(33 downto 0) := (others => '0');
signal s694 : std_logic_vector(33 downto 0) := (others => '0');
signal s695 : std_logic_vector(33 downto 0) := (others => '0');
signal s696 : std_logic_vector(33 downto 0) := (others => '0');
signal s697 : std_logic_vector(33 downto 0) := (others => '0');
signal s698 : std_logic_vector(33 downto 0) := (others => '0');
signal s699 : std_logic_vector(33 downto 0) := (others => '0');
signal s700 : std_logic_vector(33 downto 0) := (others => '0');
signal s701 : std_logic_vector(33 downto 0) := (others => '0');
signal s702 : std_logic_vector(33 downto 0) := (others => '0');
signal s703 : std_logic_vector(33 downto 0) := (others => '0');
signal s704 : std_logic_vector(33 downto 0) := (others => '0');
signal s705 : std_logic_vector(33 downto 0) := (others => '0');
signal s706 : std_logic_vector(33 downto 0) := (others => '0');
signal s707 : std_logic_vector(33 downto 0) := (others => '0');
signal s708 : std_logic_vector(33 downto 0) := (others => '0');
signal s709 : std_logic_vector(33 downto 0) := (others => '0');
signal s710 : std_logic_vector(33 downto 0) := (others => '0');
signal s711 : std_logic_vector(33 downto 0) := (others => '0');
signal s712 : std_logic_vector(33 downto 0) := (others => '0');
signal s713 : std_logic_vector(33 downto 0) := (others => '0');
signal s714 : std_logic_vector(33 downto 0) := (others => '0');
signal s715 : std_logic_vector(33 downto 0) := (others => '0');
signal s716 : std_logic_vector(33 downto 0) := (others => '0');
signal s717 : std_logic_vector(33 downto 0) := (others => '0');
signal s718 : std_logic_vector(33 downto 0) := (others => '0');
signal s719 : std_logic_vector(33 downto 0) := (others => '0');
signal s720 : std_logic_vector(33 downto 0) := (others => '0');
signal s721 : std_logic_vector(33 downto 0) := (others => '0');
signal s722 : std_logic_vector(33 downto 0) := (others => '0');
signal s723 : std_logic_vector(33 downto 0) := (others => '0');
signal s724 : std_logic_vector(33 downto 0) := (others => '0');
signal s725 : std_logic_vector(33 downto 0) := (others => '0');
signal s726 : std_logic_vector(33 downto 0) := (others => '0');
signal s727 : std_logic_vector(33 downto 0) := (others => '0');
signal s728 : std_logic_vector(33 downto 0) := (others => '0');
signal s729 : std_logic_vector(33 downto 0) := (others => '0');
signal s730 : std_logic_vector(33 downto 0) := (others => '0');
signal s731 : std_logic_vector(33 downto 0) := (others => '0');
signal s732 : std_logic_vector(33 downto 0) := (others => '0');
signal s733 : std_logic_vector(33 downto 0) := (others => '0');
signal s734 : std_logic_vector(33 downto 0) := (others => '0');
signal s735 : std_logic_vector(33 downto 0) := (others => '0');
signal s736 : std_logic_vector(33 downto 0) := (others => '0');
signal s737 : std_logic_vector(33 downto 0) := (others => '0');
signal s738 : std_logic_vector(33 downto 0) := (others => '0');
signal s739 : std_logic_vector(33 downto 0) := (others => '0');
signal s740 : std_logic_vector(33 downto 0) := (others => '0');
signal s741 : std_logic_vector(33 downto 0) := (others => '0');
signal s742 : std_logic_vector(33 downto 0) := (others => '0');
signal s743 : std_logic_vector(33 downto 0) := (others => '0');
signal s744 : std_logic_vector(33 downto 0) := (others => '0');
signal s745 : std_logic_vector(33 downto 0) := (others => '0');
signal s746 : std_logic_vector(33 downto 0) := (others => '0');
signal s747 : std_logic_vector(33 downto 0) := (others => '0');
signal s748 : std_logic_vector(33 downto 0) := (others => '0');
signal s749 : std_logic_vector(33 downto 0) := (others => '0');
signal s750 : std_logic_vector(33 downto 0) := (others => '0');
signal s751 : std_logic_vector(33 downto 0) := (others => '0');
signal s752 : std_logic_vector(33 downto 0) := (others => '0');
signal s753 : std_logic_vector(33 downto 0) := (others => '0');
signal s754 : std_logic_vector(33 downto 0) := (others => '0');
signal s755 : std_logic_vector(33 downto 0) := (others => '0');
signal s756 : std_logic_vector(33 downto 0) := (others => '0');
signal s757 : std_logic_vector(33 downto 0) := (others => '0');
signal s758 : std_logic_vector(33 downto 0) := (others => '0');
signal s759 : std_logic_vector(33 downto 0) := (others => '0');
signal s760 : std_logic_vector(33 downto 0) := (others => '0');
signal s761 : std_logic_vector(33 downto 0) := (others => '0');
signal s762 : std_logic_vector(33 downto 0) := (others => '0');
signal s763 : std_logic_vector(33 downto 0) := (others => '0');
signal s764 : std_logic_vector(33 downto 0) := (others => '0');
signal s765 : std_logic_vector(33 downto 0) := (others => '0');
signal s766 : std_logic_vector(33 downto 0) := (others => '0');
signal s767 : std_logic_vector(33 downto 0) := (others => '0');
signal s768 : std_logic_vector(33 downto 0) := (others => '0');
signal s769 : std_logic_vector(33 downto 0) := (others => '0');
signal s770 : std_logic_vector(33 downto 0) := (others => '0');
signal s771 : std_logic_vector(33 downto 0) := (others => '0');
signal s772 : std_logic_vector(33 downto 0) := (others => '0');
signal s773 : std_logic_vector(33 downto 0) := (others => '0');
signal s774 : std_logic_vector(33 downto 0) := (others => '0');
signal s775 : std_logic_vector(33 downto 0) := (others => '0');
signal s776 : std_logic_vector(33 downto 0) := (others => '0');
signal s777 : std_logic_vector(33 downto 0) := (others => '0');
signal s778 : std_logic_vector(33 downto 0) := (others => '0');
signal s779 : std_logic_vector(33 downto 0) := (others => '0');
signal s780 : std_logic_vector(33 downto 0) := (others => '0');
signal s781 : std_logic_vector(33 downto 0) := (others => '0');
signal s782 : std_logic_vector(33 downto 0) := (others => '0');
signal s783 : std_logic_vector(33 downto 0) := (others => '0');
signal s784 : std_logic_vector(33 downto 0) := (others => '0');
signal s785 : std_logic_vector(33 downto 0) := (others => '0');
signal s786 : std_logic_vector(33 downto 0) := (others => '0');
signal s787 : std_logic_vector(33 downto 0) := (others => '0');
signal s788 : std_logic_vector(33 downto 0) := (others => '0');
signal s789 : std_logic_vector(33 downto 0) := (others => '0');
signal s790 : std_logic_vector(33 downto 0) := (others => '0');
signal s791 : std_logic_vector(33 downto 0) := (others => '0');
signal s792 : std_logic_vector(33 downto 0) := (others => '0');
signal s793 : std_logic_vector(33 downto 0) := (others => '0');
signal s794 : std_logic_vector(33 downto 0) := (others => '0');
signal s795 : std_logic_vector(33 downto 0) := (others => '0');
signal s796 : std_logic_vector(33 downto 0) := (others => '0');
signal s797 : std_logic_vector(33 downto 0) := (others => '0');
signal s798 : std_logic_vector(33 downto 0) := (others => '0');
signal s799 : std_logic_vector(33 downto 0) := (others => '0');
signal s800 : std_logic_vector(33 downto 0) := (others => '0');
signal s801 : std_logic_vector(33 downto 0) := (others => '0');
signal s802 : std_logic_vector(33 downto 0) := (others => '0');
signal s803 : std_logic_vector(33 downto 0) := (others => '0');
signal s804 : std_logic_vector(33 downto 0) := (others => '0');
signal s805 : std_logic_vector(33 downto 0) := (others => '0');
signal s806 : std_logic_vector(33 downto 0) := (others => '0');
signal s807 : std_logic_vector(33 downto 0) := (others => '0');
signal s808 : std_logic_vector(33 downto 0) := (others => '0');
signal s809 : std_logic_vector(33 downto 0) := (others => '0');
signal s810 : std_logic_vector(33 downto 0) := (others => '0');
signal s811 : std_logic_vector(33 downto 0) := (others => '0');
signal s812 : std_logic_vector(33 downto 0) := (others => '0');
signal s813 : std_logic_vector(33 downto 0) := (others => '0');
signal s814 : std_logic_vector(33 downto 0) := (others => '0');
signal s815 : std_logic_vector(33 downto 0) := (others => '0');
signal s816 : std_logic_vector(33 downto 0) := (others => '0');
signal s817 : std_logic_vector(33 downto 0) := (others => '0');
signal s818 : std_logic_vector(33 downto 0) := (others => '0');
signal s819 : std_logic_vector(33 downto 0) := (others => '0');
signal s820 : std_logic_vector(33 downto 0) := (others => '0');
signal s821 : std_logic_vector(33 downto 0) := (others => '0');
signal s822 : std_logic_vector(33 downto 0) := (others => '0');
signal s823 : std_logic_vector(33 downto 0) := (others => '0');
signal s824 : std_logic_vector(33 downto 0) := (others => '0');
signal s825 : std_logic_vector(33 downto 0) := (others => '0');
signal s826 : std_logic_vector(33 downto 0) := (others => '0');
signal s827 : std_logic_vector(33 downto 0) := (others => '0');
signal s828 : std_logic_vector(33 downto 0) := (others => '0');
signal s829 : std_logic_vector(33 downto 0) := (others => '0');
signal s830 : std_logic_vector(33 downto 0) := (others => '0');
signal s831 : std_logic_vector(33 downto 0) := (others => '0');
signal s832 : std_logic_vector(33 downto 0) := (others => '0');
signal s833 : std_logic_vector(33 downto 0) := (others => '0');
signal s834 : std_logic_vector(33 downto 0) := (others => '0');
signal s835 : std_logic_vector(33 downto 0) := (others => '0');
signal s836 : std_logic_vector(33 downto 0) := (others => '0');
signal s837 : std_logic_vector(33 downto 0) := (others => '0');
signal s838 : std_logic_vector(33 downto 0) := (others => '0');
signal s839 : std_logic_vector(33 downto 0) := (others => '0');
signal s840 : std_logic_vector(33 downto 0) := (others => '0');
signal s841 : std_logic_vector(33 downto 0) := (others => '0');
signal s842 : std_logic_vector(33 downto 0) := (others => '0');
signal s843 : std_logic_vector(33 downto 0) := (others => '0');
signal s844 : std_logic_vector(33 downto 0) := (others => '0');
signal s845 : std_logic_vector(33 downto 0) := (others => '0');
signal s846 : std_logic_vector(33 downto 0) := (others => '0');
signal s847 : std_logic_vector(33 downto 0) := (others => '0');
signal s848 : std_logic_vector(33 downto 0) := (others => '0');
signal s849 : std_logic_vector(33 downto 0) := (others => '0');
signal s850 : std_logic_vector(33 downto 0) := (others => '0');
signal s851 : std_logic_vector(33 downto 0) := (others => '0');
signal s852 : std_logic_vector(33 downto 0) := (others => '0');
signal s853 : std_logic_vector(33 downto 0) := (others => '0');
signal s854 : std_logic_vector(33 downto 0) := (others => '0');
signal s855 : std_logic_vector(33 downto 0) := (others => '0');
signal s856 : std_logic_vector(33 downto 0) := (others => '0');
signal s857 : std_logic_vector(33 downto 0) := (others => '0');
signal s858 : std_logic_vector(33 downto 0) := (others => '0');
signal s859 : std_logic_vector(33 downto 0) := (others => '0');
signal s860 : std_logic_vector(33 downto 0) := (others => '0');
signal s861 : std_logic_vector(33 downto 0) := (others => '0');
signal s862 : std_logic_vector(33 downto 0) := (others => '0');
signal s863 : std_logic_vector(33 downto 0) := (others => '0');
signal s864 : std_logic_vector(33 downto 0) := (others => '0');
signal s865 : std_logic_vector(33 downto 0) := (others => '0');
signal s866 : std_logic_vector(33 downto 0) := (others => '0');
signal s867 : std_logic_vector(33 downto 0) := (others => '0');
signal s868 : std_logic_vector(33 downto 0) := (others => '0');
signal s869 : std_logic_vector(33 downto 0) := (others => '0');
signal s870 : std_logic_vector(33 downto 0) := (others => '0');
signal s871 : std_logic_vector(33 downto 0) := (others => '0');
signal s872 : std_logic_vector(33 downto 0) := (others => '0');
signal s873 : std_logic_vector(33 downto 0) := (others => '0');
signal s874 : std_logic_vector(33 downto 0) := (others => '0');
signal s875 : std_logic_vector(33 downto 0) := (others => '0');
signal s876 : std_logic_vector(33 downto 0) := (others => '0');
signal s877 : std_logic_vector(33 downto 0) := (others => '0');
signal s878 : std_logic_vector(33 downto 0) := (others => '0');
signal s879 : std_logic_vector(33 downto 0) := (others => '0');
signal s880 : std_logic_vector(33 downto 0) := (others => '0');
signal s881 : std_logic_vector(33 downto 0) := (others => '0');
signal s882 : std_logic_vector(33 downto 0) := (others => '0');
signal s883 : std_logic_vector(33 downto 0) := (others => '0');
signal s884 : std_logic_vector(33 downto 0) := (others => '0');
signal s885 : std_logic_vector(33 downto 0) := (others => '0');
signal s886 : std_logic_vector(33 downto 0) := (others => '0');
signal s887 : std_logic_vector(33 downto 0) := (others => '0');
signal s888 : std_logic_vector(33 downto 0) := (others => '0');
signal s889 : std_logic_vector(33 downto 0) := (others => '0');
signal s890 : std_logic_vector(33 downto 0) := (others => '0');
signal s891 : std_logic_vector(33 downto 0) := (others => '0');
signal s892 : std_logic_vector(33 downto 0) := (others => '0');
signal s893 : std_logic_vector(33 downto 0) := (others => '0');
signal s894 : std_logic_vector(33 downto 0) := (others => '0');
signal s895 : std_logic_vector(33 downto 0) := (others => '0');
signal s896 : std_logic_vector(33 downto 0) := (others => '0');
signal s897 : std_logic_vector(33 downto 0) := (others => '0');
signal s898 : std_logic_vector(33 downto 0) := (others => '0');
signal s899 : std_logic_vector(33 downto 0) := (others => '0');
signal s900 : std_logic_vector(33 downto 0) := (others => '0');
signal s901 : std_logic_vector(33 downto 0) := (others => '0');
signal s902 : std_logic_vector(33 downto 0) := (others => '0');
signal s903 : std_logic_vector(33 downto 0) := (others => '0');
signal s904 : std_logic_vector(33 downto 0) := (others => '0');
signal s905 : std_logic_vector(33 downto 0) := (others => '0');
signal s906 : std_logic_vector(33 downto 0) := (others => '0');
signal s907 : std_logic_vector(33 downto 0) := (others => '0');
signal s908 : std_logic_vector(33 downto 0) := (others => '0');
signal s909 : std_logic_vector(33 downto 0) := (others => '0');
signal s910 : std_logic_vector(33 downto 0) := (others => '0');
signal s911 : std_logic_vector(33 downto 0) := (others => '0');
signal s912 : std_logic_vector(33 downto 0) := (others => '0');
signal s913 : std_logic_vector(33 downto 0) := (others => '0');
signal s914 : std_logic_vector(33 downto 0) := (others => '0');
signal s915 : std_logic_vector(33 downto 0) := (others => '0');
signal s916 : std_logic_vector(33 downto 0) := (others => '0');
signal s917 : std_logic_vector(33 downto 0) := (others => '0');
signal s918 : std_logic_vector(33 downto 0) := (others => '0');
signal s919 : std_logic_vector(33 downto 0) := (others => '0');
signal s920 : std_logic_vector(33 downto 0) := (others => '0');
signal s921 : std_logic_vector(33 downto 0) := (others => '0');
signal s922 : std_logic_vector(33 downto 0) := (others => '0');
signal s923 : std_logic_vector(33 downto 0) := (others => '0');
signal s924 : std_logic_vector(33 downto 0) := (others => '0');
signal s925 : std_logic_vector(33 downto 0) := (others => '0');
signal s926 : std_logic_vector(33 downto 0) := (others => '0');
signal s927 : std_logic_vector(33 downto 0) := (others => '0');
signal s928 : std_logic_vector(33 downto 0) := (others => '0');
signal s929 : std_logic_vector(33 downto 0) := (others => '0');
signal s930 : std_logic_vector(33 downto 0) := (others => '0');
signal s931 : std_logic_vector(33 downto 0) := (others => '0');
signal s932 : std_logic_vector(33 downto 0) := (others => '0');
signal s933 : std_logic_vector(33 downto 0) := (others => '0');
signal s934 : std_logic_vector(33 downto 0) := (others => '0');
signal s935 : std_logic_vector(33 downto 0) := (others => '0');
signal s936 : std_logic_vector(33 downto 0) := (others => '0');
signal s937 : std_logic_vector(33 downto 0) := (others => '0');
signal s938 : std_logic_vector(33 downto 0) := (others => '0');
signal s939 : std_logic_vector(33 downto 0) := (others => '0');
signal s940 : std_logic_vector(33 downto 0) := (others => '0');
signal s941 : std_logic_vector(33 downto 0) := (others => '0');
signal s942 : std_logic_vector(33 downto 0) := (others => '0');
signal s943 : std_logic_vector(33 downto 0) := (others => '0');
signal s944 : std_logic_vector(33 downto 0) := (others => '0');
signal s945 : std_logic_vector(33 downto 0) := (others => '0');
signal s946 : std_logic_vector(33 downto 0) := (others => '0');
signal s947 : std_logic_vector(33 downto 0) := (others => '0');
signal s948 : std_logic_vector(33 downto 0) := (others => '0');
signal s949 : std_logic_vector(33 downto 0) := (others => '0');
signal s950 : std_logic_vector(33 downto 0) := (others => '0');
signal s951 : std_logic_vector(33 downto 0) := (others => '0');
signal s952 : std_logic_vector(33 downto 0) := (others => '0');
signal s953 : std_logic_vector(33 downto 0) := (others => '0');
signal s954 : std_logic_vector(33 downto 0) := (others => '0');
signal s955 : std_logic_vector(33 downto 0) := (others => '0');
signal s956 : std_logic_vector(33 downto 0) := (others => '0');
signal s957 : std_logic_vector(33 downto 0) := (others => '0');
signal s958 : std_logic_vector(33 downto 0) := (others => '0');
signal s959 : std_logic_vector(33 downto 0) := (others => '0');
signal s960 : std_logic_vector(33 downto 0) := (others => '0');
signal s961 : std_logic_vector(33 downto 0) := (others => '0');
signal s962 : std_logic_vector(33 downto 0) := (others => '0');
signal s963 : std_logic_vector(33 downto 0) := (others => '0');
signal s964 : std_logic_vector(33 downto 0) := (others => '0');
signal s965 : std_logic_vector(33 downto 0) := (others => '0');
signal s966 : std_logic_vector(33 downto 0) := (others => '0');
signal s967 : std_logic_vector(33 downto 0) := (others => '0');
signal s968 : std_logic_vector(33 downto 0) := (others => '0');
signal s969 : std_logic_vector(33 downto 0) := (others => '0');
signal s970 : std_logic_vector(33 downto 0) := (others => '0');
signal s971 : std_logic_vector(33 downto 0) := (others => '0');
signal s972 : std_logic_vector(33 downto 0) := (others => '0');
signal s973 : std_logic_vector(33 downto 0) := (others => '0');
signal s974 : std_logic_vector(33 downto 0) := (others => '0');
signal s975 : std_logic_vector(33 downto 0) := (others => '0');
signal s976 : std_logic_vector(33 downto 0) := (others => '0');
signal s977 : std_logic_vector(33 downto 0) := (others => '0');
signal s978 : std_logic_vector(33 downto 0) := (others => '0');
signal s979 : std_logic_vector(33 downto 0) := (others => '0');
signal s980 : std_logic_vector(33 downto 0) := (others => '0');
signal s981 : std_logic_vector(33 downto 0) := (others => '0');
signal s982 : std_logic_vector(33 downto 0) := (others => '0');
signal s983 : std_logic_vector(33 downto 0) := (others => '0');
signal s984 : std_logic_vector(33 downto 0) := (others => '0');
signal s985 : std_logic_vector(33 downto 0) := (others => '0');
signal s986 : std_logic_vector(33 downto 0) := (others => '0');
signal s987 : std_logic_vector(33 downto 0) := (others => '0');
signal s988 : std_logic_vector(33 downto 0) := (others => '0');
signal s989 : std_logic_vector(33 downto 0) := (others => '0');
signal s990 : std_logic_vector(33 downto 0) := (others => '0');
signal s991 : std_logic_vector(33 downto 0) := (others => '0');
signal s992 : std_logic_vector(33 downto 0) := (others => '0');
signal s993 : std_logic_vector(33 downto 0) := (others => '0');
signal s994 : std_logic_vector(33 downto 0) := (others => '0');
signal s995 : std_logic_vector(33 downto 0) := (others => '0');
signal s996 : std_logic_vector(33 downto 0) := (others => '0');
signal s997 : std_logic_vector(33 downto 0) := (others => '0');
signal s998 : std_logic_vector(33 downto 0) := (others => '0');
signal s999 : std_logic_vector(33 downto 0) := (others => '0');
signal s1000 : std_logic_vector(33 downto 0) := (others => '0');
signal s1001 : std_logic_vector(33 downto 0) := (others => '0');
signal s1002 : std_logic_vector(33 downto 0) := (others => '0');
signal s1003 : std_logic_vector(33 downto 0) := (others => '0');
signal s1004 : std_logic_vector(33 downto 0) := (others => '0');
signal s1005 : std_logic_vector(33 downto 0) := (others => '0');
signal s1006 : std_logic_vector(33 downto 0) := (others => '0');
signal s1007 : std_logic_vector(33 downto 0) := (others => '0');
signal s1008 : std_logic_vector(33 downto 0) := (others => '0');
signal s1009 : std_logic_vector(33 downto 0) := (others => '0');
signal s1010 : std_logic_vector(33 downto 0) := (others => '0');
signal s1011 : std_logic_vector(33 downto 0) := (others => '0');
signal s1012 : std_logic_vector(33 downto 0) := (others => '0');
signal s1013 : std_logic_vector(33 downto 0) := (others => '0');
signal s1014 : std_logic_vector(33 downto 0) := (others => '0');
signal s1015 : std_logic_vector(33 downto 0) := (others => '0');
signal s1016 : std_logic_vector(33 downto 0) := (others => '0');
signal s1017 : std_logic_vector(33 downto 0) := (others => '0');
signal s1018 : std_logic_vector(33 downto 0) := (others => '0');
signal s1019 : std_logic_vector(33 downto 0) := (others => '0');
signal s1020 : std_logic_vector(33 downto 0) := (others => '0');
signal s1021 : std_logic_vector(33 downto 0) := (others => '0');
signal s1022 : std_logic_vector(33 downto 0) := (others => '0');
signal s1023 : std_logic_vector(33 downto 0) := (others => '0');
signal s1024 : std_logic_vector(33 downto 0) := (others => '0');
signal s1025 : std_logic_vector(33 downto 0) := (others => '0');
signal s1026 : std_logic_vector(33 downto 0) := (others => '0');
signal s1027 : std_logic_vector(33 downto 0) := (others => '0');
signal s1028 : std_logic_vector(33 downto 0) := (others => '0');
signal s1029 : std_logic_vector(33 downto 0) := (others => '0');
signal s1030 : std_logic_vector(33 downto 0) := (others => '0');
signal s1031 : std_logic_vector(33 downto 0) := (others => '0');
signal s1032 : std_logic_vector(33 downto 0) := (others => '0');
signal s1033 : std_logic_vector(33 downto 0) := (others => '0');
signal s1034 : std_logic_vector(33 downto 0) := (others => '0');
signal s1035 : std_logic_vector(33 downto 0) := (others => '0');
signal s1036 : std_logic_vector(33 downto 0) := (others => '0');
signal s1037 : std_logic_vector(33 downto 0) := (others => '0');
signal s1038 : std_logic_vector(33 downto 0) := (others => '0');
signal s1039 : std_logic_vector(33 downto 0) := (others => '0');
signal s1040 : std_logic_vector(33 downto 0) := (others => '0');
signal s1041 : std_logic_vector(33 downto 0) := (others => '0');
signal s1042 : std_logic_vector(33 downto 0) := (others => '0');
signal s1043 : std_logic_vector(33 downto 0) := (others => '0');
signal s1044 : std_logic_vector(33 downto 0) := (others => '0');
signal s1045 : std_logic_vector(33 downto 0) := (others => '0');
signal s1046 : std_logic_vector(33 downto 0) := (others => '0');
signal s1047 : std_logic_vector(33 downto 0) := (others => '0');
signal s1048 : std_logic_vector(33 downto 0) := (others => '0');
signal s1049 : std_logic_vector(33 downto 0) := (others => '0');
signal s1050 : std_logic_vector(33 downto 0) := (others => '0');
signal s1051 : std_logic_vector(33 downto 0) := (others => '0');
signal s1052 : std_logic_vector(33 downto 0) := (others => '0');
signal s1053 : std_logic_vector(33 downto 0) := (others => '0');
signal s1054 : std_logic_vector(33 downto 0) := (others => '0');
signal s1055 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
      s558 <= "0000000000000000000000000000000000";
      s559 <= "0000000000000000000000000000000000";
      s560 <= "0000000000000000000000000000000000";
      s561 <= "0000000000000000000000000000000000";
      s562 <= "0000000000000000000000000000000000";
      s563 <= "0000000000000000000000000000000000";
      s564 <= "0000000000000000000000000000000000";
      s565 <= "0000000000000000000000000000000000";
      s566 <= "0000000000000000000000000000000000";
      s567 <= "0000000000000000000000000000000000";
      s568 <= "0000000000000000000000000000000000";
      s569 <= "0000000000000000000000000000000000";
      s570 <= "0000000000000000000000000000000000";
      s571 <= "0000000000000000000000000000000000";
      s572 <= "0000000000000000000000000000000000";
      s573 <= "0000000000000000000000000000000000";
      s574 <= "0000000000000000000000000000000000";
      s575 <= "0000000000000000000000000000000000";
      s576 <= "0000000000000000000000000000000000";
      s577 <= "0000000000000000000000000000000000";
      s578 <= "0000000000000000000000000000000000";
      s579 <= "0000000000000000000000000000000000";
      s580 <= "0000000000000000000000000000000000";
      s581 <= "0000000000000000000000000000000000";
      s582 <= "0000000000000000000000000000000000";
      s583 <= "0000000000000000000000000000000000";
      s584 <= "0000000000000000000000000000000000";
      s585 <= "0000000000000000000000000000000000";
      s586 <= "0000000000000000000000000000000000";
      s587 <= "0000000000000000000000000000000000";
      s588 <= "0000000000000000000000000000000000";
      s589 <= "0000000000000000000000000000000000";
      s590 <= "0000000000000000000000000000000000";
      s591 <= "0000000000000000000000000000000000";
      s592 <= "0000000000000000000000000000000000";
      s593 <= "0000000000000000000000000000000000";
      s594 <= "0000000000000000000000000000000000";
      s595 <= "0000000000000000000000000000000000";
      s596 <= "0000000000000000000000000000000000";
      s597 <= "0000000000000000000000000000000000";
      s598 <= "0000000000000000000000000000000000";
      s599 <= "0000000000000000000000000000000000";
      s600 <= "0000000000000000000000000000000000";
      s601 <= "0000000000000000000000000000000000";
      s602 <= "0000000000000000000000000000000000";
      s603 <= "0000000000000000000000000000000000";
      s604 <= "0000000000000000000000000000000000";
      s605 <= "0000000000000000000000000000000000";
      s606 <= "0000000000000000000000000000000000";
      s607 <= "0000000000000000000000000000000000";
      s608 <= "0000000000000000000000000000000000";
      s609 <= "0000000000000000000000000000000000";
      s610 <= "0000000000000000000000000000000000";
      s611 <= "0000000000000000000000000000000000";
      s612 <= "0000000000000000000000000000000000";
      s613 <= "0000000000000000000000000000000000";
      s614 <= "0000000000000000000000000000000000";
      s615 <= "0000000000000000000000000000000000";
      s616 <= "0000000000000000000000000000000000";
      s617 <= "0000000000000000000000000000000000";
      s618 <= "0000000000000000000000000000000000";
      s619 <= "0000000000000000000000000000000000";
      s620 <= "0000000000000000000000000000000000";
      s621 <= "0000000000000000000000000000000000";
      s622 <= "0000000000000000000000000000000000";
      s623 <= "0000000000000000000000000000000000";
      s624 <= "0000000000000000000000000000000000";
      s625 <= "0000000000000000000000000000000000";
      s626 <= "0000000000000000000000000000000000";
      s627 <= "0000000000000000000000000000000000";
      s628 <= "0000000000000000000000000000000000";
      s629 <= "0000000000000000000000000000000000";
      s630 <= "0000000000000000000000000000000000";
      s631 <= "0000000000000000000000000000000000";
      s632 <= "0000000000000000000000000000000000";
      s633 <= "0000000000000000000000000000000000";
      s634 <= "0000000000000000000000000000000000";
      s635 <= "0000000000000000000000000000000000";
      s636 <= "0000000000000000000000000000000000";
      s637 <= "0000000000000000000000000000000000";
      s638 <= "0000000000000000000000000000000000";
      s639 <= "0000000000000000000000000000000000";
      s640 <= "0000000000000000000000000000000000";
      s641 <= "0000000000000000000000000000000000";
      s642 <= "0000000000000000000000000000000000";
      s643 <= "0000000000000000000000000000000000";
      s644 <= "0000000000000000000000000000000000";
      s645 <= "0000000000000000000000000000000000";
      s646 <= "0000000000000000000000000000000000";
      s647 <= "0000000000000000000000000000000000";
      s648 <= "0000000000000000000000000000000000";
      s649 <= "0000000000000000000000000000000000";
      s650 <= "0000000000000000000000000000000000";
      s651 <= "0000000000000000000000000000000000";
      s652 <= "0000000000000000000000000000000000";
      s653 <= "0000000000000000000000000000000000";
      s654 <= "0000000000000000000000000000000000";
      s655 <= "0000000000000000000000000000000000";
      s656 <= "0000000000000000000000000000000000";
      s657 <= "0000000000000000000000000000000000";
      s658 <= "0000000000000000000000000000000000";
      s659 <= "0000000000000000000000000000000000";
      s660 <= "0000000000000000000000000000000000";
      s661 <= "0000000000000000000000000000000000";
      s662 <= "0000000000000000000000000000000000";
      s663 <= "0000000000000000000000000000000000";
      s664 <= "0000000000000000000000000000000000";
      s665 <= "0000000000000000000000000000000000";
      s666 <= "0000000000000000000000000000000000";
      s667 <= "0000000000000000000000000000000000";
      s668 <= "0000000000000000000000000000000000";
      s669 <= "0000000000000000000000000000000000";
      s670 <= "0000000000000000000000000000000000";
      s671 <= "0000000000000000000000000000000000";
      s672 <= "0000000000000000000000000000000000";
      s673 <= "0000000000000000000000000000000000";
      s674 <= "0000000000000000000000000000000000";
      s675 <= "0000000000000000000000000000000000";
      s676 <= "0000000000000000000000000000000000";
      s677 <= "0000000000000000000000000000000000";
      s678 <= "0000000000000000000000000000000000";
      s679 <= "0000000000000000000000000000000000";
      s680 <= "0000000000000000000000000000000000";
      s681 <= "0000000000000000000000000000000000";
      s682 <= "0000000000000000000000000000000000";
      s683 <= "0000000000000000000000000000000000";
      s684 <= "0000000000000000000000000000000000";
      s685 <= "0000000000000000000000000000000000";
      s686 <= "0000000000000000000000000000000000";
      s687 <= "0000000000000000000000000000000000";
      s688 <= "0000000000000000000000000000000000";
      s689 <= "0000000000000000000000000000000000";
      s690 <= "0000000000000000000000000000000000";
      s691 <= "0000000000000000000000000000000000";
      s692 <= "0000000000000000000000000000000000";
      s693 <= "0000000000000000000000000000000000";
      s694 <= "0000000000000000000000000000000000";
      s695 <= "0000000000000000000000000000000000";
      s696 <= "0000000000000000000000000000000000";
      s697 <= "0000000000000000000000000000000000";
      s698 <= "0000000000000000000000000000000000";
      s699 <= "0000000000000000000000000000000000";
      s700 <= "0000000000000000000000000000000000";
      s701 <= "0000000000000000000000000000000000";
      s702 <= "0000000000000000000000000000000000";
      s703 <= "0000000000000000000000000000000000";
      s704 <= "0000000000000000000000000000000000";
      s705 <= "0000000000000000000000000000000000";
      s706 <= "0000000000000000000000000000000000";
      s707 <= "0000000000000000000000000000000000";
      s708 <= "0000000000000000000000000000000000";
      s709 <= "0000000000000000000000000000000000";
      s710 <= "0000000000000000000000000000000000";
      s711 <= "0000000000000000000000000000000000";
      s712 <= "0000000000000000000000000000000000";
      s713 <= "0000000000000000000000000000000000";
      s714 <= "0000000000000000000000000000000000";
      s715 <= "0000000000000000000000000000000000";
      s716 <= "0000000000000000000000000000000000";
      s717 <= "0000000000000000000000000000000000";
      s718 <= "0000000000000000000000000000000000";
      s719 <= "0000000000000000000000000000000000";
      s720 <= "0000000000000000000000000000000000";
      s721 <= "0000000000000000000000000000000000";
      s722 <= "0000000000000000000000000000000000";
      s723 <= "0000000000000000000000000000000000";
      s724 <= "0000000000000000000000000000000000";
      s725 <= "0000000000000000000000000000000000";
      s726 <= "0000000000000000000000000000000000";
      s727 <= "0000000000000000000000000000000000";
      s728 <= "0000000000000000000000000000000000";
      s729 <= "0000000000000000000000000000000000";
      s730 <= "0000000000000000000000000000000000";
      s731 <= "0000000000000000000000000000000000";
      s732 <= "0000000000000000000000000000000000";
      s733 <= "0000000000000000000000000000000000";
      s734 <= "0000000000000000000000000000000000";
      s735 <= "0000000000000000000000000000000000";
      s736 <= "0000000000000000000000000000000000";
      s737 <= "0000000000000000000000000000000000";
      s738 <= "0000000000000000000000000000000000";
      s739 <= "0000000000000000000000000000000000";
      s740 <= "0000000000000000000000000000000000";
      s741 <= "0000000000000000000000000000000000";
      s742 <= "0000000000000000000000000000000000";
      s743 <= "0000000000000000000000000000000000";
      s744 <= "0000000000000000000000000000000000";
      s745 <= "0000000000000000000000000000000000";
      s746 <= "0000000000000000000000000000000000";
      s747 <= "0000000000000000000000000000000000";
      s748 <= "0000000000000000000000000000000000";
      s749 <= "0000000000000000000000000000000000";
      s750 <= "0000000000000000000000000000000000";
      s751 <= "0000000000000000000000000000000000";
      s752 <= "0000000000000000000000000000000000";
      s753 <= "0000000000000000000000000000000000";
      s754 <= "0000000000000000000000000000000000";
      s755 <= "0000000000000000000000000000000000";
      s756 <= "0000000000000000000000000000000000";
      s757 <= "0000000000000000000000000000000000";
      s758 <= "0000000000000000000000000000000000";
      s759 <= "0000000000000000000000000000000000";
      s760 <= "0000000000000000000000000000000000";
      s761 <= "0000000000000000000000000000000000";
      s762 <= "0000000000000000000000000000000000";
      s763 <= "0000000000000000000000000000000000";
      s764 <= "0000000000000000000000000000000000";
      s765 <= "0000000000000000000000000000000000";
      s766 <= "0000000000000000000000000000000000";
      s767 <= "0000000000000000000000000000000000";
      s768 <= "0000000000000000000000000000000000";
      s769 <= "0000000000000000000000000000000000";
      s770 <= "0000000000000000000000000000000000";
      s771 <= "0000000000000000000000000000000000";
      s772 <= "0000000000000000000000000000000000";
      s773 <= "0000000000000000000000000000000000";
      s774 <= "0000000000000000000000000000000000";
      s775 <= "0000000000000000000000000000000000";
      s776 <= "0000000000000000000000000000000000";
      s777 <= "0000000000000000000000000000000000";
      s778 <= "0000000000000000000000000000000000";
      s779 <= "0000000000000000000000000000000000";
      s780 <= "0000000000000000000000000000000000";
      s781 <= "0000000000000000000000000000000000";
      s782 <= "0000000000000000000000000000000000";
      s783 <= "0000000000000000000000000000000000";
      s784 <= "0000000000000000000000000000000000";
      s785 <= "0000000000000000000000000000000000";
      s786 <= "0000000000000000000000000000000000";
      s787 <= "0000000000000000000000000000000000";
      s788 <= "0000000000000000000000000000000000";
      s789 <= "0000000000000000000000000000000000";
      s790 <= "0000000000000000000000000000000000";
      s791 <= "0000000000000000000000000000000000";
      s792 <= "0000000000000000000000000000000000";
      s793 <= "0000000000000000000000000000000000";
      s794 <= "0000000000000000000000000000000000";
      s795 <= "0000000000000000000000000000000000";
      s796 <= "0000000000000000000000000000000000";
      s797 <= "0000000000000000000000000000000000";
      s798 <= "0000000000000000000000000000000000";
      s799 <= "0000000000000000000000000000000000";
      s800 <= "0000000000000000000000000000000000";
      s801 <= "0000000000000000000000000000000000";
      s802 <= "0000000000000000000000000000000000";
      s803 <= "0000000000000000000000000000000000";
      s804 <= "0000000000000000000000000000000000";
      s805 <= "0000000000000000000000000000000000";
      s806 <= "0000000000000000000000000000000000";
      s807 <= "0000000000000000000000000000000000";
      s808 <= "0000000000000000000000000000000000";
      s809 <= "0000000000000000000000000000000000";
      s810 <= "0000000000000000000000000000000000";
      s811 <= "0000000000000000000000000000000000";
      s812 <= "0000000000000000000000000000000000";
      s813 <= "0000000000000000000000000000000000";
      s814 <= "0000000000000000000000000000000000";
      s815 <= "0000000000000000000000000000000000";
      s816 <= "0000000000000000000000000000000000";
      s817 <= "0000000000000000000000000000000000";
      s818 <= "0000000000000000000000000000000000";
      s819 <= "0000000000000000000000000000000000";
      s820 <= "0000000000000000000000000000000000";
      s821 <= "0000000000000000000000000000000000";
      s822 <= "0000000000000000000000000000000000";
      s823 <= "0000000000000000000000000000000000";
      s824 <= "0000000000000000000000000000000000";
      s825 <= "0000000000000000000000000000000000";
      s826 <= "0000000000000000000000000000000000";
      s827 <= "0000000000000000000000000000000000";
      s828 <= "0000000000000000000000000000000000";
      s829 <= "0000000000000000000000000000000000";
      s830 <= "0000000000000000000000000000000000";
      s831 <= "0000000000000000000000000000000000";
      s832 <= "0000000000000000000000000000000000";
      s833 <= "0000000000000000000000000000000000";
      s834 <= "0000000000000000000000000000000000";
      s835 <= "0000000000000000000000000000000000";
      s836 <= "0000000000000000000000000000000000";
      s837 <= "0000000000000000000000000000000000";
      s838 <= "0000000000000000000000000000000000";
      s839 <= "0000000000000000000000000000000000";
      s840 <= "0000000000000000000000000000000000";
      s841 <= "0000000000000000000000000000000000";
      s842 <= "0000000000000000000000000000000000";
      s843 <= "0000000000000000000000000000000000";
      s844 <= "0000000000000000000000000000000000";
      s845 <= "0000000000000000000000000000000000";
      s846 <= "0000000000000000000000000000000000";
      s847 <= "0000000000000000000000000000000000";
      s848 <= "0000000000000000000000000000000000";
      s849 <= "0000000000000000000000000000000000";
      s850 <= "0000000000000000000000000000000000";
      s851 <= "0000000000000000000000000000000000";
      s852 <= "0000000000000000000000000000000000";
      s853 <= "0000000000000000000000000000000000";
      s854 <= "0000000000000000000000000000000000";
      s855 <= "0000000000000000000000000000000000";
      s856 <= "0000000000000000000000000000000000";
      s857 <= "0000000000000000000000000000000000";
      s858 <= "0000000000000000000000000000000000";
      s859 <= "0000000000000000000000000000000000";
      s860 <= "0000000000000000000000000000000000";
      s861 <= "0000000000000000000000000000000000";
      s862 <= "0000000000000000000000000000000000";
      s863 <= "0000000000000000000000000000000000";
      s864 <= "0000000000000000000000000000000000";
      s865 <= "0000000000000000000000000000000000";
      s866 <= "0000000000000000000000000000000000";
      s867 <= "0000000000000000000000000000000000";
      s868 <= "0000000000000000000000000000000000";
      s869 <= "0000000000000000000000000000000000";
      s870 <= "0000000000000000000000000000000000";
      s871 <= "0000000000000000000000000000000000";
      s872 <= "0000000000000000000000000000000000";
      s873 <= "0000000000000000000000000000000000";
      s874 <= "0000000000000000000000000000000000";
      s875 <= "0000000000000000000000000000000000";
      s876 <= "0000000000000000000000000000000000";
      s877 <= "0000000000000000000000000000000000";
      s878 <= "0000000000000000000000000000000000";
      s879 <= "0000000000000000000000000000000000";
      s880 <= "0000000000000000000000000000000000";
      s881 <= "0000000000000000000000000000000000";
      s882 <= "0000000000000000000000000000000000";
      s883 <= "0000000000000000000000000000000000";
      s884 <= "0000000000000000000000000000000000";
      s885 <= "0000000000000000000000000000000000";
      s886 <= "0000000000000000000000000000000000";
      s887 <= "0000000000000000000000000000000000";
      s888 <= "0000000000000000000000000000000000";
      s889 <= "0000000000000000000000000000000000";
      s890 <= "0000000000000000000000000000000000";
      s891 <= "0000000000000000000000000000000000";
      s892 <= "0000000000000000000000000000000000";
      s893 <= "0000000000000000000000000000000000";
      s894 <= "0000000000000000000000000000000000";
      s895 <= "0000000000000000000000000000000000";
      s896 <= "0000000000000000000000000000000000";
      s897 <= "0000000000000000000000000000000000";
      s898 <= "0000000000000000000000000000000000";
      s899 <= "0000000000000000000000000000000000";
      s900 <= "0000000000000000000000000000000000";
      s901 <= "0000000000000000000000000000000000";
      s902 <= "0000000000000000000000000000000000";
      s903 <= "0000000000000000000000000000000000";
      s904 <= "0000000000000000000000000000000000";
      s905 <= "0000000000000000000000000000000000";
      s906 <= "0000000000000000000000000000000000";
      s907 <= "0000000000000000000000000000000000";
      s908 <= "0000000000000000000000000000000000";
      s909 <= "0000000000000000000000000000000000";
      s910 <= "0000000000000000000000000000000000";
      s911 <= "0000000000000000000000000000000000";
      s912 <= "0000000000000000000000000000000000";
      s913 <= "0000000000000000000000000000000000";
      s914 <= "0000000000000000000000000000000000";
      s915 <= "0000000000000000000000000000000000";
      s916 <= "0000000000000000000000000000000000";
      s917 <= "0000000000000000000000000000000000";
      s918 <= "0000000000000000000000000000000000";
      s919 <= "0000000000000000000000000000000000";
      s920 <= "0000000000000000000000000000000000";
      s921 <= "0000000000000000000000000000000000";
      s922 <= "0000000000000000000000000000000000";
      s923 <= "0000000000000000000000000000000000";
      s924 <= "0000000000000000000000000000000000";
      s925 <= "0000000000000000000000000000000000";
      s926 <= "0000000000000000000000000000000000";
      s927 <= "0000000000000000000000000000000000";
      s928 <= "0000000000000000000000000000000000";
      s929 <= "0000000000000000000000000000000000";
      s930 <= "0000000000000000000000000000000000";
      s931 <= "0000000000000000000000000000000000";
      s932 <= "0000000000000000000000000000000000";
      s933 <= "0000000000000000000000000000000000";
      s934 <= "0000000000000000000000000000000000";
      s935 <= "0000000000000000000000000000000000";
      s936 <= "0000000000000000000000000000000000";
      s937 <= "0000000000000000000000000000000000";
      s938 <= "0000000000000000000000000000000000";
      s939 <= "0000000000000000000000000000000000";
      s940 <= "0000000000000000000000000000000000";
      s941 <= "0000000000000000000000000000000000";
      s942 <= "0000000000000000000000000000000000";
      s943 <= "0000000000000000000000000000000000";
      s944 <= "0000000000000000000000000000000000";
      s945 <= "0000000000000000000000000000000000";
      s946 <= "0000000000000000000000000000000000";
      s947 <= "0000000000000000000000000000000000";
      s948 <= "0000000000000000000000000000000000";
      s949 <= "0000000000000000000000000000000000";
      s950 <= "0000000000000000000000000000000000";
      s951 <= "0000000000000000000000000000000000";
      s952 <= "0000000000000000000000000000000000";
      s953 <= "0000000000000000000000000000000000";
      s954 <= "0000000000000000000000000000000000";
      s955 <= "0000000000000000000000000000000000";
      s956 <= "0000000000000000000000000000000000";
      s957 <= "0000000000000000000000000000000000";
      s958 <= "0000000000000000000000000000000000";
      s959 <= "0000000000000000000000000000000000";
      s960 <= "0000000000000000000000000000000000";
      s961 <= "0000000000000000000000000000000000";
      s962 <= "0000000000000000000000000000000000";
      s963 <= "0000000000000000000000000000000000";
      s964 <= "0000000000000000000000000000000000";
      s965 <= "0000000000000000000000000000000000";
      s966 <= "0000000000000000000000000000000000";
      s967 <= "0000000000000000000000000000000000";
      s968 <= "0000000000000000000000000000000000";
      s969 <= "0000000000000000000000000000000000";
      s970 <= "0000000000000000000000000000000000";
      s971 <= "0000000000000000000000000000000000";
      s972 <= "0000000000000000000000000000000000";
      s973 <= "0000000000000000000000000000000000";
      s974 <= "0000000000000000000000000000000000";
      s975 <= "0000000000000000000000000000000000";
      s976 <= "0000000000000000000000000000000000";
      s977 <= "0000000000000000000000000000000000";
      s978 <= "0000000000000000000000000000000000";
      s979 <= "0000000000000000000000000000000000";
      s980 <= "0000000000000000000000000000000000";
      s981 <= "0000000000000000000000000000000000";
      s982 <= "0000000000000000000000000000000000";
      s983 <= "0000000000000000000000000000000000";
      s984 <= "0000000000000000000000000000000000";
      s985 <= "0000000000000000000000000000000000";
      s986 <= "0000000000000000000000000000000000";
      s987 <= "0000000000000000000000000000000000";
      s988 <= "0000000000000000000000000000000000";
      s989 <= "0000000000000000000000000000000000";
      s990 <= "0000000000000000000000000000000000";
      s991 <= "0000000000000000000000000000000000";
      s992 <= "0000000000000000000000000000000000";
      s993 <= "0000000000000000000000000000000000";
      s994 <= "0000000000000000000000000000000000";
      s995 <= "0000000000000000000000000000000000";
      s996 <= "0000000000000000000000000000000000";
      s997 <= "0000000000000000000000000000000000";
      s998 <= "0000000000000000000000000000000000";
      s999 <= "0000000000000000000000000000000000";
      s1000 <= "0000000000000000000000000000000000";
      s1001 <= "0000000000000000000000000000000000";
      s1002 <= "0000000000000000000000000000000000";
      s1003 <= "0000000000000000000000000000000000";
      s1004 <= "0000000000000000000000000000000000";
      s1005 <= "0000000000000000000000000000000000";
      s1006 <= "0000000000000000000000000000000000";
      s1007 <= "0000000000000000000000000000000000";
      s1008 <= "0000000000000000000000000000000000";
      s1009 <= "0000000000000000000000000000000000";
      s1010 <= "0000000000000000000000000000000000";
      s1011 <= "0000000000000000000000000000000000";
      s1012 <= "0000000000000000000000000000000000";
      s1013 <= "0000000000000000000000000000000000";
      s1014 <= "0000000000000000000000000000000000";
      s1015 <= "0000000000000000000000000000000000";
      s1016 <= "0000000000000000000000000000000000";
      s1017 <= "0000000000000000000000000000000000";
      s1018 <= "0000000000000000000000000000000000";
      s1019 <= "0000000000000000000000000000000000";
      s1020 <= "0000000000000000000000000000000000";
      s1021 <= "0000000000000000000000000000000000";
      s1022 <= "0000000000000000000000000000000000";
      s1023 <= "0000000000000000000000000000000000";
      s1024 <= "0000000000000000000000000000000000";
      s1025 <= "0000000000000000000000000000000000";
      s1026 <= "0000000000000000000000000000000000";
      s1027 <= "0000000000000000000000000000000000";
      s1028 <= "0000000000000000000000000000000000";
      s1029 <= "0000000000000000000000000000000000";
      s1030 <= "0000000000000000000000000000000000";
      s1031 <= "0000000000000000000000000000000000";
      s1032 <= "0000000000000000000000000000000000";
      s1033 <= "0000000000000000000000000000000000";
      s1034 <= "0000000000000000000000000000000000";
      s1035 <= "0000000000000000000000000000000000";
      s1036 <= "0000000000000000000000000000000000";
      s1037 <= "0000000000000000000000000000000000";
      s1038 <= "0000000000000000000000000000000000";
      s1039 <= "0000000000000000000000000000000000";
      s1040 <= "0000000000000000000000000000000000";
      s1041 <= "0000000000000000000000000000000000";
      s1042 <= "0000000000000000000000000000000000";
      s1043 <= "0000000000000000000000000000000000";
      s1044 <= "0000000000000000000000000000000000";
      s1045 <= "0000000000000000000000000000000000";
      s1046 <= "0000000000000000000000000000000000";
      s1047 <= "0000000000000000000000000000000000";
      s1048 <= "0000000000000000000000000000000000";
      s1049 <= "0000000000000000000000000000000000";
      s1050 <= "0000000000000000000000000000000000";
      s1051 <= "0000000000000000000000000000000000";
      s1052 <= "0000000000000000000000000000000000";
      s1053 <= "0000000000000000000000000000000000";
      s1054 <= "0000000000000000000000000000000000";
      s1055 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      s558 <= s557;
      s559 <= s558;
      s560 <= s559;
      s561 <= s560;
      s562 <= s561;
      s563 <= s562;
      s564 <= s563;
      s565 <= s564;
      s566 <= s565;
      s567 <= s566;
      s568 <= s567;
      s569 <= s568;
      s570 <= s569;
      s571 <= s570;
      s572 <= s571;
      s573 <= s572;
      s574 <= s573;
      s575 <= s574;
      s576 <= s575;
      s577 <= s576;
      s578 <= s577;
      s579 <= s578;
      s580 <= s579;
      s581 <= s580;
      s582 <= s581;
      s583 <= s582;
      s584 <= s583;
      s585 <= s584;
      s586 <= s585;
      s587 <= s586;
      s588 <= s587;
      s589 <= s588;
      s590 <= s589;
      s591 <= s590;
      s592 <= s591;
      s593 <= s592;
      s594 <= s593;
      s595 <= s594;
      s596 <= s595;
      s597 <= s596;
      s598 <= s597;
      s599 <= s598;
      s600 <= s599;
      s601 <= s600;
      s602 <= s601;
      s603 <= s602;
      s604 <= s603;
      s605 <= s604;
      s606 <= s605;
      s607 <= s606;
      s608 <= s607;
      s609 <= s608;
      s610 <= s609;
      s611 <= s610;
      s612 <= s611;
      s613 <= s612;
      s614 <= s613;
      s615 <= s614;
      s616 <= s615;
      s617 <= s616;
      s618 <= s617;
      s619 <= s618;
      s620 <= s619;
      s621 <= s620;
      s622 <= s621;
      s623 <= s622;
      s624 <= s623;
      s625 <= s624;
      s626 <= s625;
      s627 <= s626;
      s628 <= s627;
      s629 <= s628;
      s630 <= s629;
      s631 <= s630;
      s632 <= s631;
      s633 <= s632;
      s634 <= s633;
      s635 <= s634;
      s636 <= s635;
      s637 <= s636;
      s638 <= s637;
      s639 <= s638;
      s640 <= s639;
      s641 <= s640;
      s642 <= s641;
      s643 <= s642;
      s644 <= s643;
      s645 <= s644;
      s646 <= s645;
      s647 <= s646;
      s648 <= s647;
      s649 <= s648;
      s650 <= s649;
      s651 <= s650;
      s652 <= s651;
      s653 <= s652;
      s654 <= s653;
      s655 <= s654;
      s656 <= s655;
      s657 <= s656;
      s658 <= s657;
      s659 <= s658;
      s660 <= s659;
      s661 <= s660;
      s662 <= s661;
      s663 <= s662;
      s664 <= s663;
      s665 <= s664;
      s666 <= s665;
      s667 <= s666;
      s668 <= s667;
      s669 <= s668;
      s670 <= s669;
      s671 <= s670;
      s672 <= s671;
      s673 <= s672;
      s674 <= s673;
      s675 <= s674;
      s676 <= s675;
      s677 <= s676;
      s678 <= s677;
      s679 <= s678;
      s680 <= s679;
      s681 <= s680;
      s682 <= s681;
      s683 <= s682;
      s684 <= s683;
      s685 <= s684;
      s686 <= s685;
      s687 <= s686;
      s688 <= s687;
      s689 <= s688;
      s690 <= s689;
      s691 <= s690;
      s692 <= s691;
      s693 <= s692;
      s694 <= s693;
      s695 <= s694;
      s696 <= s695;
      s697 <= s696;
      s698 <= s697;
      s699 <= s698;
      s700 <= s699;
      s701 <= s700;
      s702 <= s701;
      s703 <= s702;
      s704 <= s703;
      s705 <= s704;
      s706 <= s705;
      s707 <= s706;
      s708 <= s707;
      s709 <= s708;
      s710 <= s709;
      s711 <= s710;
      s712 <= s711;
      s713 <= s712;
      s714 <= s713;
      s715 <= s714;
      s716 <= s715;
      s717 <= s716;
      s718 <= s717;
      s719 <= s718;
      s720 <= s719;
      s721 <= s720;
      s722 <= s721;
      s723 <= s722;
      s724 <= s723;
      s725 <= s724;
      s726 <= s725;
      s727 <= s726;
      s728 <= s727;
      s729 <= s728;
      s730 <= s729;
      s731 <= s730;
      s732 <= s731;
      s733 <= s732;
      s734 <= s733;
      s735 <= s734;
      s736 <= s735;
      s737 <= s736;
      s738 <= s737;
      s739 <= s738;
      s740 <= s739;
      s741 <= s740;
      s742 <= s741;
      s743 <= s742;
      s744 <= s743;
      s745 <= s744;
      s746 <= s745;
      s747 <= s746;
      s748 <= s747;
      s749 <= s748;
      s750 <= s749;
      s751 <= s750;
      s752 <= s751;
      s753 <= s752;
      s754 <= s753;
      s755 <= s754;
      s756 <= s755;
      s757 <= s756;
      s758 <= s757;
      s759 <= s758;
      s760 <= s759;
      s761 <= s760;
      s762 <= s761;
      s763 <= s762;
      s764 <= s763;
      s765 <= s764;
      s766 <= s765;
      s767 <= s766;
      s768 <= s767;
      s769 <= s768;
      s770 <= s769;
      s771 <= s770;
      s772 <= s771;
      s773 <= s772;
      s774 <= s773;
      s775 <= s774;
      s776 <= s775;
      s777 <= s776;
      s778 <= s777;
      s779 <= s778;
      s780 <= s779;
      s781 <= s780;
      s782 <= s781;
      s783 <= s782;
      s784 <= s783;
      s785 <= s784;
      s786 <= s785;
      s787 <= s786;
      s788 <= s787;
      s789 <= s788;
      s790 <= s789;
      s791 <= s790;
      s792 <= s791;
      s793 <= s792;
      s794 <= s793;
      s795 <= s794;
      s796 <= s795;
      s797 <= s796;
      s798 <= s797;
      s799 <= s798;
      s800 <= s799;
      s801 <= s800;
      s802 <= s801;
      s803 <= s802;
      s804 <= s803;
      s805 <= s804;
      s806 <= s805;
      s807 <= s806;
      s808 <= s807;
      s809 <= s808;
      s810 <= s809;
      s811 <= s810;
      s812 <= s811;
      s813 <= s812;
      s814 <= s813;
      s815 <= s814;
      s816 <= s815;
      s817 <= s816;
      s818 <= s817;
      s819 <= s818;
      s820 <= s819;
      s821 <= s820;
      s822 <= s821;
      s823 <= s822;
      s824 <= s823;
      s825 <= s824;
      s826 <= s825;
      s827 <= s826;
      s828 <= s827;
      s829 <= s828;
      s830 <= s829;
      s831 <= s830;
      s832 <= s831;
      s833 <= s832;
      s834 <= s833;
      s835 <= s834;
      s836 <= s835;
      s837 <= s836;
      s838 <= s837;
      s839 <= s838;
      s840 <= s839;
      s841 <= s840;
      s842 <= s841;
      s843 <= s842;
      s844 <= s843;
      s845 <= s844;
      s846 <= s845;
      s847 <= s846;
      s848 <= s847;
      s849 <= s848;
      s850 <= s849;
      s851 <= s850;
      s852 <= s851;
      s853 <= s852;
      s854 <= s853;
      s855 <= s854;
      s856 <= s855;
      s857 <= s856;
      s858 <= s857;
      s859 <= s858;
      s860 <= s859;
      s861 <= s860;
      s862 <= s861;
      s863 <= s862;
      s864 <= s863;
      s865 <= s864;
      s866 <= s865;
      s867 <= s866;
      s868 <= s867;
      s869 <= s868;
      s870 <= s869;
      s871 <= s870;
      s872 <= s871;
      s873 <= s872;
      s874 <= s873;
      s875 <= s874;
      s876 <= s875;
      s877 <= s876;
      s878 <= s877;
      s879 <= s878;
      s880 <= s879;
      s881 <= s880;
      s882 <= s881;
      s883 <= s882;
      s884 <= s883;
      s885 <= s884;
      s886 <= s885;
      s887 <= s886;
      s888 <= s887;
      s889 <= s888;
      s890 <= s889;
      s891 <= s890;
      s892 <= s891;
      s893 <= s892;
      s894 <= s893;
      s895 <= s894;
      s896 <= s895;
      s897 <= s896;
      s898 <= s897;
      s899 <= s898;
      s900 <= s899;
      s901 <= s900;
      s902 <= s901;
      s903 <= s902;
      s904 <= s903;
      s905 <= s904;
      s906 <= s905;
      s907 <= s906;
      s908 <= s907;
      s909 <= s908;
      s910 <= s909;
      s911 <= s910;
      s912 <= s911;
      s913 <= s912;
      s914 <= s913;
      s915 <= s914;
      s916 <= s915;
      s917 <= s916;
      s918 <= s917;
      s919 <= s918;
      s920 <= s919;
      s921 <= s920;
      s922 <= s921;
      s923 <= s922;
      s924 <= s923;
      s925 <= s924;
      s926 <= s925;
      s927 <= s926;
      s928 <= s927;
      s929 <= s928;
      s930 <= s929;
      s931 <= s930;
      s932 <= s931;
      s933 <= s932;
      s934 <= s933;
      s935 <= s934;
      s936 <= s935;
      s937 <= s936;
      s938 <= s937;
      s939 <= s938;
      s940 <= s939;
      s941 <= s940;
      s942 <= s941;
      s943 <= s942;
      s944 <= s943;
      s945 <= s944;
      s946 <= s945;
      s947 <= s946;
      s948 <= s947;
      s949 <= s948;
      s950 <= s949;
      s951 <= s950;
      s952 <= s951;
      s953 <= s952;
      s954 <= s953;
      s955 <= s954;
      s956 <= s955;
      s957 <= s956;
      s958 <= s957;
      s959 <= s958;
      s960 <= s959;
      s961 <= s960;
      s962 <= s961;
      s963 <= s962;
      s964 <= s963;
      s965 <= s964;
      s966 <= s965;
      s967 <= s966;
      s968 <= s967;
      s969 <= s968;
      s970 <= s969;
      s971 <= s970;
      s972 <= s971;
      s973 <= s972;
      s974 <= s973;
      s975 <= s974;
      s976 <= s975;
      s977 <= s976;
      s978 <= s977;
      s979 <= s978;
      s980 <= s979;
      s981 <= s980;
      s982 <= s981;
      s983 <= s982;
      s984 <= s983;
      s985 <= s984;
      s986 <= s985;
      s987 <= s986;
      s988 <= s987;
      s989 <= s988;
      s990 <= s989;
      s991 <= s990;
      s992 <= s991;
      s993 <= s992;
      s994 <= s993;
      s995 <= s994;
      s996 <= s995;
      s997 <= s996;
      s998 <= s997;
      s999 <= s998;
      s1000 <= s999;
      s1001 <= s1000;
      s1002 <= s1001;
      s1003 <= s1002;
      s1004 <= s1003;
      s1005 <= s1004;
      s1006 <= s1005;
      s1007 <= s1006;
      s1008 <= s1007;
      s1009 <= s1008;
      s1010 <= s1009;
      s1011 <= s1010;
      s1012 <= s1011;
      s1013 <= s1012;
      s1014 <= s1013;
      s1015 <= s1014;
      s1016 <= s1015;
      s1017 <= s1016;
      s1018 <= s1017;
      s1019 <= s1018;
      s1020 <= s1019;
      s1021 <= s1020;
      s1022 <= s1021;
      s1023 <= s1022;
      s1024 <= s1023;
      s1025 <= s1024;
      s1026 <= s1025;
      s1027 <= s1026;
      s1028 <= s1027;
      s1029 <= s1028;
      s1030 <= s1029;
      s1031 <= s1030;
      s1032 <= s1031;
      s1033 <= s1032;
      s1034 <= s1033;
      s1035 <= s1034;
      s1036 <= s1035;
      s1037 <= s1036;
      s1038 <= s1037;
      s1039 <= s1038;
      s1040 <= s1039;
      s1041 <= s1040;
      s1042 <= s1041;
      s1043 <= s1042;
      s1044 <= s1043;
      s1045 <= s1044;
      s1046 <= s1045;
      s1047 <= s1046;
      s1048 <= s1047;
      s1049 <= s1048;
      s1050 <= s1049;
      s1051 <= s1050;
      s1052 <= s1051;
      s1053 <= s1052;
      s1054 <= s1053;
      s1055 <= s1054;
      Y <= s1055;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_146_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 146 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_146_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_146_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      Y <= s145;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_239_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 239 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_239_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_239_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      Y <= s238;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_294_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 294 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_294_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_294_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      Y <= s293;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_359_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 359 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_359_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_359_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      Y <= s358;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_442_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 442 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_442_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_442_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      Y <= s441;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_499_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 499 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_499_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_499_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      Y <= s498;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_555_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 555 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_555_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_555_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      Y <= s554;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_625_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 625 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_625_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_625_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
signal s165 : std_logic_vector(33 downto 0) := (others => '0');
signal s166 : std_logic_vector(33 downto 0) := (others => '0');
signal s167 : std_logic_vector(33 downto 0) := (others => '0');
signal s168 : std_logic_vector(33 downto 0) := (others => '0');
signal s169 : std_logic_vector(33 downto 0) := (others => '0');
signal s170 : std_logic_vector(33 downto 0) := (others => '0');
signal s171 : std_logic_vector(33 downto 0) := (others => '0');
signal s172 : std_logic_vector(33 downto 0) := (others => '0');
signal s173 : std_logic_vector(33 downto 0) := (others => '0');
signal s174 : std_logic_vector(33 downto 0) := (others => '0');
signal s175 : std_logic_vector(33 downto 0) := (others => '0');
signal s176 : std_logic_vector(33 downto 0) := (others => '0');
signal s177 : std_logic_vector(33 downto 0) := (others => '0');
signal s178 : std_logic_vector(33 downto 0) := (others => '0');
signal s179 : std_logic_vector(33 downto 0) := (others => '0');
signal s180 : std_logic_vector(33 downto 0) := (others => '0');
signal s181 : std_logic_vector(33 downto 0) := (others => '0');
signal s182 : std_logic_vector(33 downto 0) := (others => '0');
signal s183 : std_logic_vector(33 downto 0) := (others => '0');
signal s184 : std_logic_vector(33 downto 0) := (others => '0');
signal s185 : std_logic_vector(33 downto 0) := (others => '0');
signal s186 : std_logic_vector(33 downto 0) := (others => '0');
signal s187 : std_logic_vector(33 downto 0) := (others => '0');
signal s188 : std_logic_vector(33 downto 0) := (others => '0');
signal s189 : std_logic_vector(33 downto 0) := (others => '0');
signal s190 : std_logic_vector(33 downto 0) := (others => '0');
signal s191 : std_logic_vector(33 downto 0) := (others => '0');
signal s192 : std_logic_vector(33 downto 0) := (others => '0');
signal s193 : std_logic_vector(33 downto 0) := (others => '0');
signal s194 : std_logic_vector(33 downto 0) := (others => '0');
signal s195 : std_logic_vector(33 downto 0) := (others => '0');
signal s196 : std_logic_vector(33 downto 0) := (others => '0');
signal s197 : std_logic_vector(33 downto 0) := (others => '0');
signal s198 : std_logic_vector(33 downto 0) := (others => '0');
signal s199 : std_logic_vector(33 downto 0) := (others => '0');
signal s200 : std_logic_vector(33 downto 0) := (others => '0');
signal s201 : std_logic_vector(33 downto 0) := (others => '0');
signal s202 : std_logic_vector(33 downto 0) := (others => '0');
signal s203 : std_logic_vector(33 downto 0) := (others => '0');
signal s204 : std_logic_vector(33 downto 0) := (others => '0');
signal s205 : std_logic_vector(33 downto 0) := (others => '0');
signal s206 : std_logic_vector(33 downto 0) := (others => '0');
signal s207 : std_logic_vector(33 downto 0) := (others => '0');
signal s208 : std_logic_vector(33 downto 0) := (others => '0');
signal s209 : std_logic_vector(33 downto 0) := (others => '0');
signal s210 : std_logic_vector(33 downto 0) := (others => '0');
signal s211 : std_logic_vector(33 downto 0) := (others => '0');
signal s212 : std_logic_vector(33 downto 0) := (others => '0');
signal s213 : std_logic_vector(33 downto 0) := (others => '0');
signal s214 : std_logic_vector(33 downto 0) := (others => '0');
signal s215 : std_logic_vector(33 downto 0) := (others => '0');
signal s216 : std_logic_vector(33 downto 0) := (others => '0');
signal s217 : std_logic_vector(33 downto 0) := (others => '0');
signal s218 : std_logic_vector(33 downto 0) := (others => '0');
signal s219 : std_logic_vector(33 downto 0) := (others => '0');
signal s220 : std_logic_vector(33 downto 0) := (others => '0');
signal s221 : std_logic_vector(33 downto 0) := (others => '0');
signal s222 : std_logic_vector(33 downto 0) := (others => '0');
signal s223 : std_logic_vector(33 downto 0) := (others => '0');
signal s224 : std_logic_vector(33 downto 0) := (others => '0');
signal s225 : std_logic_vector(33 downto 0) := (others => '0');
signal s226 : std_logic_vector(33 downto 0) := (others => '0');
signal s227 : std_logic_vector(33 downto 0) := (others => '0');
signal s228 : std_logic_vector(33 downto 0) := (others => '0');
signal s229 : std_logic_vector(33 downto 0) := (others => '0');
signal s230 : std_logic_vector(33 downto 0) := (others => '0');
signal s231 : std_logic_vector(33 downto 0) := (others => '0');
signal s232 : std_logic_vector(33 downto 0) := (others => '0');
signal s233 : std_logic_vector(33 downto 0) := (others => '0');
signal s234 : std_logic_vector(33 downto 0) := (others => '0');
signal s235 : std_logic_vector(33 downto 0) := (others => '0');
signal s236 : std_logic_vector(33 downto 0) := (others => '0');
signal s237 : std_logic_vector(33 downto 0) := (others => '0');
signal s238 : std_logic_vector(33 downto 0) := (others => '0');
signal s239 : std_logic_vector(33 downto 0) := (others => '0');
signal s240 : std_logic_vector(33 downto 0) := (others => '0');
signal s241 : std_logic_vector(33 downto 0) := (others => '0');
signal s242 : std_logic_vector(33 downto 0) := (others => '0');
signal s243 : std_logic_vector(33 downto 0) := (others => '0');
signal s244 : std_logic_vector(33 downto 0) := (others => '0');
signal s245 : std_logic_vector(33 downto 0) := (others => '0');
signal s246 : std_logic_vector(33 downto 0) := (others => '0');
signal s247 : std_logic_vector(33 downto 0) := (others => '0');
signal s248 : std_logic_vector(33 downto 0) := (others => '0');
signal s249 : std_logic_vector(33 downto 0) := (others => '0');
signal s250 : std_logic_vector(33 downto 0) := (others => '0');
signal s251 : std_logic_vector(33 downto 0) := (others => '0');
signal s252 : std_logic_vector(33 downto 0) := (others => '0');
signal s253 : std_logic_vector(33 downto 0) := (others => '0');
signal s254 : std_logic_vector(33 downto 0) := (others => '0');
signal s255 : std_logic_vector(33 downto 0) := (others => '0');
signal s256 : std_logic_vector(33 downto 0) := (others => '0');
signal s257 : std_logic_vector(33 downto 0) := (others => '0');
signal s258 : std_logic_vector(33 downto 0) := (others => '0');
signal s259 : std_logic_vector(33 downto 0) := (others => '0');
signal s260 : std_logic_vector(33 downto 0) := (others => '0');
signal s261 : std_logic_vector(33 downto 0) := (others => '0');
signal s262 : std_logic_vector(33 downto 0) := (others => '0');
signal s263 : std_logic_vector(33 downto 0) := (others => '0');
signal s264 : std_logic_vector(33 downto 0) := (others => '0');
signal s265 : std_logic_vector(33 downto 0) := (others => '0');
signal s266 : std_logic_vector(33 downto 0) := (others => '0');
signal s267 : std_logic_vector(33 downto 0) := (others => '0');
signal s268 : std_logic_vector(33 downto 0) := (others => '0');
signal s269 : std_logic_vector(33 downto 0) := (others => '0');
signal s270 : std_logic_vector(33 downto 0) := (others => '0');
signal s271 : std_logic_vector(33 downto 0) := (others => '0');
signal s272 : std_logic_vector(33 downto 0) := (others => '0');
signal s273 : std_logic_vector(33 downto 0) := (others => '0');
signal s274 : std_logic_vector(33 downto 0) := (others => '0');
signal s275 : std_logic_vector(33 downto 0) := (others => '0');
signal s276 : std_logic_vector(33 downto 0) := (others => '0');
signal s277 : std_logic_vector(33 downto 0) := (others => '0');
signal s278 : std_logic_vector(33 downto 0) := (others => '0');
signal s279 : std_logic_vector(33 downto 0) := (others => '0');
signal s280 : std_logic_vector(33 downto 0) := (others => '0');
signal s281 : std_logic_vector(33 downto 0) := (others => '0');
signal s282 : std_logic_vector(33 downto 0) := (others => '0');
signal s283 : std_logic_vector(33 downto 0) := (others => '0');
signal s284 : std_logic_vector(33 downto 0) := (others => '0');
signal s285 : std_logic_vector(33 downto 0) := (others => '0');
signal s286 : std_logic_vector(33 downto 0) := (others => '0');
signal s287 : std_logic_vector(33 downto 0) := (others => '0');
signal s288 : std_logic_vector(33 downto 0) := (others => '0');
signal s289 : std_logic_vector(33 downto 0) := (others => '0');
signal s290 : std_logic_vector(33 downto 0) := (others => '0');
signal s291 : std_logic_vector(33 downto 0) := (others => '0');
signal s292 : std_logic_vector(33 downto 0) := (others => '0');
signal s293 : std_logic_vector(33 downto 0) := (others => '0');
signal s294 : std_logic_vector(33 downto 0) := (others => '0');
signal s295 : std_logic_vector(33 downto 0) := (others => '0');
signal s296 : std_logic_vector(33 downto 0) := (others => '0');
signal s297 : std_logic_vector(33 downto 0) := (others => '0');
signal s298 : std_logic_vector(33 downto 0) := (others => '0');
signal s299 : std_logic_vector(33 downto 0) := (others => '0');
signal s300 : std_logic_vector(33 downto 0) := (others => '0');
signal s301 : std_logic_vector(33 downto 0) := (others => '0');
signal s302 : std_logic_vector(33 downto 0) := (others => '0');
signal s303 : std_logic_vector(33 downto 0) := (others => '0');
signal s304 : std_logic_vector(33 downto 0) := (others => '0');
signal s305 : std_logic_vector(33 downto 0) := (others => '0');
signal s306 : std_logic_vector(33 downto 0) := (others => '0');
signal s307 : std_logic_vector(33 downto 0) := (others => '0');
signal s308 : std_logic_vector(33 downto 0) := (others => '0');
signal s309 : std_logic_vector(33 downto 0) := (others => '0');
signal s310 : std_logic_vector(33 downto 0) := (others => '0');
signal s311 : std_logic_vector(33 downto 0) := (others => '0');
signal s312 : std_logic_vector(33 downto 0) := (others => '0');
signal s313 : std_logic_vector(33 downto 0) := (others => '0');
signal s314 : std_logic_vector(33 downto 0) := (others => '0');
signal s315 : std_logic_vector(33 downto 0) := (others => '0');
signal s316 : std_logic_vector(33 downto 0) := (others => '0');
signal s317 : std_logic_vector(33 downto 0) := (others => '0');
signal s318 : std_logic_vector(33 downto 0) := (others => '0');
signal s319 : std_logic_vector(33 downto 0) := (others => '0');
signal s320 : std_logic_vector(33 downto 0) := (others => '0');
signal s321 : std_logic_vector(33 downto 0) := (others => '0');
signal s322 : std_logic_vector(33 downto 0) := (others => '0');
signal s323 : std_logic_vector(33 downto 0) := (others => '0');
signal s324 : std_logic_vector(33 downto 0) := (others => '0');
signal s325 : std_logic_vector(33 downto 0) := (others => '0');
signal s326 : std_logic_vector(33 downto 0) := (others => '0');
signal s327 : std_logic_vector(33 downto 0) := (others => '0');
signal s328 : std_logic_vector(33 downto 0) := (others => '0');
signal s329 : std_logic_vector(33 downto 0) := (others => '0');
signal s330 : std_logic_vector(33 downto 0) := (others => '0');
signal s331 : std_logic_vector(33 downto 0) := (others => '0');
signal s332 : std_logic_vector(33 downto 0) := (others => '0');
signal s333 : std_logic_vector(33 downto 0) := (others => '0');
signal s334 : std_logic_vector(33 downto 0) := (others => '0');
signal s335 : std_logic_vector(33 downto 0) := (others => '0');
signal s336 : std_logic_vector(33 downto 0) := (others => '0');
signal s337 : std_logic_vector(33 downto 0) := (others => '0');
signal s338 : std_logic_vector(33 downto 0) := (others => '0');
signal s339 : std_logic_vector(33 downto 0) := (others => '0');
signal s340 : std_logic_vector(33 downto 0) := (others => '0');
signal s341 : std_logic_vector(33 downto 0) := (others => '0');
signal s342 : std_logic_vector(33 downto 0) := (others => '0');
signal s343 : std_logic_vector(33 downto 0) := (others => '0');
signal s344 : std_logic_vector(33 downto 0) := (others => '0');
signal s345 : std_logic_vector(33 downto 0) := (others => '0');
signal s346 : std_logic_vector(33 downto 0) := (others => '0');
signal s347 : std_logic_vector(33 downto 0) := (others => '0');
signal s348 : std_logic_vector(33 downto 0) := (others => '0');
signal s349 : std_logic_vector(33 downto 0) := (others => '0');
signal s350 : std_logic_vector(33 downto 0) := (others => '0');
signal s351 : std_logic_vector(33 downto 0) := (others => '0');
signal s352 : std_logic_vector(33 downto 0) := (others => '0');
signal s353 : std_logic_vector(33 downto 0) := (others => '0');
signal s354 : std_logic_vector(33 downto 0) := (others => '0');
signal s355 : std_logic_vector(33 downto 0) := (others => '0');
signal s356 : std_logic_vector(33 downto 0) := (others => '0');
signal s357 : std_logic_vector(33 downto 0) := (others => '0');
signal s358 : std_logic_vector(33 downto 0) := (others => '0');
signal s359 : std_logic_vector(33 downto 0) := (others => '0');
signal s360 : std_logic_vector(33 downto 0) := (others => '0');
signal s361 : std_logic_vector(33 downto 0) := (others => '0');
signal s362 : std_logic_vector(33 downto 0) := (others => '0');
signal s363 : std_logic_vector(33 downto 0) := (others => '0');
signal s364 : std_logic_vector(33 downto 0) := (others => '0');
signal s365 : std_logic_vector(33 downto 0) := (others => '0');
signal s366 : std_logic_vector(33 downto 0) := (others => '0');
signal s367 : std_logic_vector(33 downto 0) := (others => '0');
signal s368 : std_logic_vector(33 downto 0) := (others => '0');
signal s369 : std_logic_vector(33 downto 0) := (others => '0');
signal s370 : std_logic_vector(33 downto 0) := (others => '0');
signal s371 : std_logic_vector(33 downto 0) := (others => '0');
signal s372 : std_logic_vector(33 downto 0) := (others => '0');
signal s373 : std_logic_vector(33 downto 0) := (others => '0');
signal s374 : std_logic_vector(33 downto 0) := (others => '0');
signal s375 : std_logic_vector(33 downto 0) := (others => '0');
signal s376 : std_logic_vector(33 downto 0) := (others => '0');
signal s377 : std_logic_vector(33 downto 0) := (others => '0');
signal s378 : std_logic_vector(33 downto 0) := (others => '0');
signal s379 : std_logic_vector(33 downto 0) := (others => '0');
signal s380 : std_logic_vector(33 downto 0) := (others => '0');
signal s381 : std_logic_vector(33 downto 0) := (others => '0');
signal s382 : std_logic_vector(33 downto 0) := (others => '0');
signal s383 : std_logic_vector(33 downto 0) := (others => '0');
signal s384 : std_logic_vector(33 downto 0) := (others => '0');
signal s385 : std_logic_vector(33 downto 0) := (others => '0');
signal s386 : std_logic_vector(33 downto 0) := (others => '0');
signal s387 : std_logic_vector(33 downto 0) := (others => '0');
signal s388 : std_logic_vector(33 downto 0) := (others => '0');
signal s389 : std_logic_vector(33 downto 0) := (others => '0');
signal s390 : std_logic_vector(33 downto 0) := (others => '0');
signal s391 : std_logic_vector(33 downto 0) := (others => '0');
signal s392 : std_logic_vector(33 downto 0) := (others => '0');
signal s393 : std_logic_vector(33 downto 0) := (others => '0');
signal s394 : std_logic_vector(33 downto 0) := (others => '0');
signal s395 : std_logic_vector(33 downto 0) := (others => '0');
signal s396 : std_logic_vector(33 downto 0) := (others => '0');
signal s397 : std_logic_vector(33 downto 0) := (others => '0');
signal s398 : std_logic_vector(33 downto 0) := (others => '0');
signal s399 : std_logic_vector(33 downto 0) := (others => '0');
signal s400 : std_logic_vector(33 downto 0) := (others => '0');
signal s401 : std_logic_vector(33 downto 0) := (others => '0');
signal s402 : std_logic_vector(33 downto 0) := (others => '0');
signal s403 : std_logic_vector(33 downto 0) := (others => '0');
signal s404 : std_logic_vector(33 downto 0) := (others => '0');
signal s405 : std_logic_vector(33 downto 0) := (others => '0');
signal s406 : std_logic_vector(33 downto 0) := (others => '0');
signal s407 : std_logic_vector(33 downto 0) := (others => '0');
signal s408 : std_logic_vector(33 downto 0) := (others => '0');
signal s409 : std_logic_vector(33 downto 0) := (others => '0');
signal s410 : std_logic_vector(33 downto 0) := (others => '0');
signal s411 : std_logic_vector(33 downto 0) := (others => '0');
signal s412 : std_logic_vector(33 downto 0) := (others => '0');
signal s413 : std_logic_vector(33 downto 0) := (others => '0');
signal s414 : std_logic_vector(33 downto 0) := (others => '0');
signal s415 : std_logic_vector(33 downto 0) := (others => '0');
signal s416 : std_logic_vector(33 downto 0) := (others => '0');
signal s417 : std_logic_vector(33 downto 0) := (others => '0');
signal s418 : std_logic_vector(33 downto 0) := (others => '0');
signal s419 : std_logic_vector(33 downto 0) := (others => '0');
signal s420 : std_logic_vector(33 downto 0) := (others => '0');
signal s421 : std_logic_vector(33 downto 0) := (others => '0');
signal s422 : std_logic_vector(33 downto 0) := (others => '0');
signal s423 : std_logic_vector(33 downto 0) := (others => '0');
signal s424 : std_logic_vector(33 downto 0) := (others => '0');
signal s425 : std_logic_vector(33 downto 0) := (others => '0');
signal s426 : std_logic_vector(33 downto 0) := (others => '0');
signal s427 : std_logic_vector(33 downto 0) := (others => '0');
signal s428 : std_logic_vector(33 downto 0) := (others => '0');
signal s429 : std_logic_vector(33 downto 0) := (others => '0');
signal s430 : std_logic_vector(33 downto 0) := (others => '0');
signal s431 : std_logic_vector(33 downto 0) := (others => '0');
signal s432 : std_logic_vector(33 downto 0) := (others => '0');
signal s433 : std_logic_vector(33 downto 0) := (others => '0');
signal s434 : std_logic_vector(33 downto 0) := (others => '0');
signal s435 : std_logic_vector(33 downto 0) := (others => '0');
signal s436 : std_logic_vector(33 downto 0) := (others => '0');
signal s437 : std_logic_vector(33 downto 0) := (others => '0');
signal s438 : std_logic_vector(33 downto 0) := (others => '0');
signal s439 : std_logic_vector(33 downto 0) := (others => '0');
signal s440 : std_logic_vector(33 downto 0) := (others => '0');
signal s441 : std_logic_vector(33 downto 0) := (others => '0');
signal s442 : std_logic_vector(33 downto 0) := (others => '0');
signal s443 : std_logic_vector(33 downto 0) := (others => '0');
signal s444 : std_logic_vector(33 downto 0) := (others => '0');
signal s445 : std_logic_vector(33 downto 0) := (others => '0');
signal s446 : std_logic_vector(33 downto 0) := (others => '0');
signal s447 : std_logic_vector(33 downto 0) := (others => '0');
signal s448 : std_logic_vector(33 downto 0) := (others => '0');
signal s449 : std_logic_vector(33 downto 0) := (others => '0');
signal s450 : std_logic_vector(33 downto 0) := (others => '0');
signal s451 : std_logic_vector(33 downto 0) := (others => '0');
signal s452 : std_logic_vector(33 downto 0) := (others => '0');
signal s453 : std_logic_vector(33 downto 0) := (others => '0');
signal s454 : std_logic_vector(33 downto 0) := (others => '0');
signal s455 : std_logic_vector(33 downto 0) := (others => '0');
signal s456 : std_logic_vector(33 downto 0) := (others => '0');
signal s457 : std_logic_vector(33 downto 0) := (others => '0');
signal s458 : std_logic_vector(33 downto 0) := (others => '0');
signal s459 : std_logic_vector(33 downto 0) := (others => '0');
signal s460 : std_logic_vector(33 downto 0) := (others => '0');
signal s461 : std_logic_vector(33 downto 0) := (others => '0');
signal s462 : std_logic_vector(33 downto 0) := (others => '0');
signal s463 : std_logic_vector(33 downto 0) := (others => '0');
signal s464 : std_logic_vector(33 downto 0) := (others => '0');
signal s465 : std_logic_vector(33 downto 0) := (others => '0');
signal s466 : std_logic_vector(33 downto 0) := (others => '0');
signal s467 : std_logic_vector(33 downto 0) := (others => '0');
signal s468 : std_logic_vector(33 downto 0) := (others => '0');
signal s469 : std_logic_vector(33 downto 0) := (others => '0');
signal s470 : std_logic_vector(33 downto 0) := (others => '0');
signal s471 : std_logic_vector(33 downto 0) := (others => '0');
signal s472 : std_logic_vector(33 downto 0) := (others => '0');
signal s473 : std_logic_vector(33 downto 0) := (others => '0');
signal s474 : std_logic_vector(33 downto 0) := (others => '0');
signal s475 : std_logic_vector(33 downto 0) := (others => '0');
signal s476 : std_logic_vector(33 downto 0) := (others => '0');
signal s477 : std_logic_vector(33 downto 0) := (others => '0');
signal s478 : std_logic_vector(33 downto 0) := (others => '0');
signal s479 : std_logic_vector(33 downto 0) := (others => '0');
signal s480 : std_logic_vector(33 downto 0) := (others => '0');
signal s481 : std_logic_vector(33 downto 0) := (others => '0');
signal s482 : std_logic_vector(33 downto 0) := (others => '0');
signal s483 : std_logic_vector(33 downto 0) := (others => '0');
signal s484 : std_logic_vector(33 downto 0) := (others => '0');
signal s485 : std_logic_vector(33 downto 0) := (others => '0');
signal s486 : std_logic_vector(33 downto 0) := (others => '0');
signal s487 : std_logic_vector(33 downto 0) := (others => '0');
signal s488 : std_logic_vector(33 downto 0) := (others => '0');
signal s489 : std_logic_vector(33 downto 0) := (others => '0');
signal s490 : std_logic_vector(33 downto 0) := (others => '0');
signal s491 : std_logic_vector(33 downto 0) := (others => '0');
signal s492 : std_logic_vector(33 downto 0) := (others => '0');
signal s493 : std_logic_vector(33 downto 0) := (others => '0');
signal s494 : std_logic_vector(33 downto 0) := (others => '0');
signal s495 : std_logic_vector(33 downto 0) := (others => '0');
signal s496 : std_logic_vector(33 downto 0) := (others => '0');
signal s497 : std_logic_vector(33 downto 0) := (others => '0');
signal s498 : std_logic_vector(33 downto 0) := (others => '0');
signal s499 : std_logic_vector(33 downto 0) := (others => '0');
signal s500 : std_logic_vector(33 downto 0) := (others => '0');
signal s501 : std_logic_vector(33 downto 0) := (others => '0');
signal s502 : std_logic_vector(33 downto 0) := (others => '0');
signal s503 : std_logic_vector(33 downto 0) := (others => '0');
signal s504 : std_logic_vector(33 downto 0) := (others => '0');
signal s505 : std_logic_vector(33 downto 0) := (others => '0');
signal s506 : std_logic_vector(33 downto 0) := (others => '0');
signal s507 : std_logic_vector(33 downto 0) := (others => '0');
signal s508 : std_logic_vector(33 downto 0) := (others => '0');
signal s509 : std_logic_vector(33 downto 0) := (others => '0');
signal s510 : std_logic_vector(33 downto 0) := (others => '0');
signal s511 : std_logic_vector(33 downto 0) := (others => '0');
signal s512 : std_logic_vector(33 downto 0) := (others => '0');
signal s513 : std_logic_vector(33 downto 0) := (others => '0');
signal s514 : std_logic_vector(33 downto 0) := (others => '0');
signal s515 : std_logic_vector(33 downto 0) := (others => '0');
signal s516 : std_logic_vector(33 downto 0) := (others => '0');
signal s517 : std_logic_vector(33 downto 0) := (others => '0');
signal s518 : std_logic_vector(33 downto 0) := (others => '0');
signal s519 : std_logic_vector(33 downto 0) := (others => '0');
signal s520 : std_logic_vector(33 downto 0) := (others => '0');
signal s521 : std_logic_vector(33 downto 0) := (others => '0');
signal s522 : std_logic_vector(33 downto 0) := (others => '0');
signal s523 : std_logic_vector(33 downto 0) := (others => '0');
signal s524 : std_logic_vector(33 downto 0) := (others => '0');
signal s525 : std_logic_vector(33 downto 0) := (others => '0');
signal s526 : std_logic_vector(33 downto 0) := (others => '0');
signal s527 : std_logic_vector(33 downto 0) := (others => '0');
signal s528 : std_logic_vector(33 downto 0) := (others => '0');
signal s529 : std_logic_vector(33 downto 0) := (others => '0');
signal s530 : std_logic_vector(33 downto 0) := (others => '0');
signal s531 : std_logic_vector(33 downto 0) := (others => '0');
signal s532 : std_logic_vector(33 downto 0) := (others => '0');
signal s533 : std_logic_vector(33 downto 0) := (others => '0');
signal s534 : std_logic_vector(33 downto 0) := (others => '0');
signal s535 : std_logic_vector(33 downto 0) := (others => '0');
signal s536 : std_logic_vector(33 downto 0) := (others => '0');
signal s537 : std_logic_vector(33 downto 0) := (others => '0');
signal s538 : std_logic_vector(33 downto 0) := (others => '0');
signal s539 : std_logic_vector(33 downto 0) := (others => '0');
signal s540 : std_logic_vector(33 downto 0) := (others => '0');
signal s541 : std_logic_vector(33 downto 0) := (others => '0');
signal s542 : std_logic_vector(33 downto 0) := (others => '0');
signal s543 : std_logic_vector(33 downto 0) := (others => '0');
signal s544 : std_logic_vector(33 downto 0) := (others => '0');
signal s545 : std_logic_vector(33 downto 0) := (others => '0');
signal s546 : std_logic_vector(33 downto 0) := (others => '0');
signal s547 : std_logic_vector(33 downto 0) := (others => '0');
signal s548 : std_logic_vector(33 downto 0) := (others => '0');
signal s549 : std_logic_vector(33 downto 0) := (others => '0');
signal s550 : std_logic_vector(33 downto 0) := (others => '0');
signal s551 : std_logic_vector(33 downto 0) := (others => '0');
signal s552 : std_logic_vector(33 downto 0) := (others => '0');
signal s553 : std_logic_vector(33 downto 0) := (others => '0');
signal s554 : std_logic_vector(33 downto 0) := (others => '0');
signal s555 : std_logic_vector(33 downto 0) := (others => '0');
signal s556 : std_logic_vector(33 downto 0) := (others => '0');
signal s557 : std_logic_vector(33 downto 0) := (others => '0');
signal s558 : std_logic_vector(33 downto 0) := (others => '0');
signal s559 : std_logic_vector(33 downto 0) := (others => '0');
signal s560 : std_logic_vector(33 downto 0) := (others => '0');
signal s561 : std_logic_vector(33 downto 0) := (others => '0');
signal s562 : std_logic_vector(33 downto 0) := (others => '0');
signal s563 : std_logic_vector(33 downto 0) := (others => '0');
signal s564 : std_logic_vector(33 downto 0) := (others => '0');
signal s565 : std_logic_vector(33 downto 0) := (others => '0');
signal s566 : std_logic_vector(33 downto 0) := (others => '0');
signal s567 : std_logic_vector(33 downto 0) := (others => '0');
signal s568 : std_logic_vector(33 downto 0) := (others => '0');
signal s569 : std_logic_vector(33 downto 0) := (others => '0');
signal s570 : std_logic_vector(33 downto 0) := (others => '0');
signal s571 : std_logic_vector(33 downto 0) := (others => '0');
signal s572 : std_logic_vector(33 downto 0) := (others => '0');
signal s573 : std_logic_vector(33 downto 0) := (others => '0');
signal s574 : std_logic_vector(33 downto 0) := (others => '0');
signal s575 : std_logic_vector(33 downto 0) := (others => '0');
signal s576 : std_logic_vector(33 downto 0) := (others => '0');
signal s577 : std_logic_vector(33 downto 0) := (others => '0');
signal s578 : std_logic_vector(33 downto 0) := (others => '0');
signal s579 : std_logic_vector(33 downto 0) := (others => '0');
signal s580 : std_logic_vector(33 downto 0) := (others => '0');
signal s581 : std_logic_vector(33 downto 0) := (others => '0');
signal s582 : std_logic_vector(33 downto 0) := (others => '0');
signal s583 : std_logic_vector(33 downto 0) := (others => '0');
signal s584 : std_logic_vector(33 downto 0) := (others => '0');
signal s585 : std_logic_vector(33 downto 0) := (others => '0');
signal s586 : std_logic_vector(33 downto 0) := (others => '0');
signal s587 : std_logic_vector(33 downto 0) := (others => '0');
signal s588 : std_logic_vector(33 downto 0) := (others => '0');
signal s589 : std_logic_vector(33 downto 0) := (others => '0');
signal s590 : std_logic_vector(33 downto 0) := (others => '0');
signal s591 : std_logic_vector(33 downto 0) := (others => '0');
signal s592 : std_logic_vector(33 downto 0) := (others => '0');
signal s593 : std_logic_vector(33 downto 0) := (others => '0');
signal s594 : std_logic_vector(33 downto 0) := (others => '0');
signal s595 : std_logic_vector(33 downto 0) := (others => '0');
signal s596 : std_logic_vector(33 downto 0) := (others => '0');
signal s597 : std_logic_vector(33 downto 0) := (others => '0');
signal s598 : std_logic_vector(33 downto 0) := (others => '0');
signal s599 : std_logic_vector(33 downto 0) := (others => '0');
signal s600 : std_logic_vector(33 downto 0) := (others => '0');
signal s601 : std_logic_vector(33 downto 0) := (others => '0');
signal s602 : std_logic_vector(33 downto 0) := (others => '0');
signal s603 : std_logic_vector(33 downto 0) := (others => '0');
signal s604 : std_logic_vector(33 downto 0) := (others => '0');
signal s605 : std_logic_vector(33 downto 0) := (others => '0');
signal s606 : std_logic_vector(33 downto 0) := (others => '0');
signal s607 : std_logic_vector(33 downto 0) := (others => '0');
signal s608 : std_logic_vector(33 downto 0) := (others => '0');
signal s609 : std_logic_vector(33 downto 0) := (others => '0');
signal s610 : std_logic_vector(33 downto 0) := (others => '0');
signal s611 : std_logic_vector(33 downto 0) := (others => '0');
signal s612 : std_logic_vector(33 downto 0) := (others => '0');
signal s613 : std_logic_vector(33 downto 0) := (others => '0');
signal s614 : std_logic_vector(33 downto 0) := (others => '0');
signal s615 : std_logic_vector(33 downto 0) := (others => '0');
signal s616 : std_logic_vector(33 downto 0) := (others => '0');
signal s617 : std_logic_vector(33 downto 0) := (others => '0');
signal s618 : std_logic_vector(33 downto 0) := (others => '0');
signal s619 : std_logic_vector(33 downto 0) := (others => '0');
signal s620 : std_logic_vector(33 downto 0) := (others => '0');
signal s621 : std_logic_vector(33 downto 0) := (others => '0');
signal s622 : std_logic_vector(33 downto 0) := (others => '0');
signal s623 : std_logic_vector(33 downto 0) := (others => '0');
signal s624 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
      s165 <= "0000000000000000000000000000000000";
      s166 <= "0000000000000000000000000000000000";
      s167 <= "0000000000000000000000000000000000";
      s168 <= "0000000000000000000000000000000000";
      s169 <= "0000000000000000000000000000000000";
      s170 <= "0000000000000000000000000000000000";
      s171 <= "0000000000000000000000000000000000";
      s172 <= "0000000000000000000000000000000000";
      s173 <= "0000000000000000000000000000000000";
      s174 <= "0000000000000000000000000000000000";
      s175 <= "0000000000000000000000000000000000";
      s176 <= "0000000000000000000000000000000000";
      s177 <= "0000000000000000000000000000000000";
      s178 <= "0000000000000000000000000000000000";
      s179 <= "0000000000000000000000000000000000";
      s180 <= "0000000000000000000000000000000000";
      s181 <= "0000000000000000000000000000000000";
      s182 <= "0000000000000000000000000000000000";
      s183 <= "0000000000000000000000000000000000";
      s184 <= "0000000000000000000000000000000000";
      s185 <= "0000000000000000000000000000000000";
      s186 <= "0000000000000000000000000000000000";
      s187 <= "0000000000000000000000000000000000";
      s188 <= "0000000000000000000000000000000000";
      s189 <= "0000000000000000000000000000000000";
      s190 <= "0000000000000000000000000000000000";
      s191 <= "0000000000000000000000000000000000";
      s192 <= "0000000000000000000000000000000000";
      s193 <= "0000000000000000000000000000000000";
      s194 <= "0000000000000000000000000000000000";
      s195 <= "0000000000000000000000000000000000";
      s196 <= "0000000000000000000000000000000000";
      s197 <= "0000000000000000000000000000000000";
      s198 <= "0000000000000000000000000000000000";
      s199 <= "0000000000000000000000000000000000";
      s200 <= "0000000000000000000000000000000000";
      s201 <= "0000000000000000000000000000000000";
      s202 <= "0000000000000000000000000000000000";
      s203 <= "0000000000000000000000000000000000";
      s204 <= "0000000000000000000000000000000000";
      s205 <= "0000000000000000000000000000000000";
      s206 <= "0000000000000000000000000000000000";
      s207 <= "0000000000000000000000000000000000";
      s208 <= "0000000000000000000000000000000000";
      s209 <= "0000000000000000000000000000000000";
      s210 <= "0000000000000000000000000000000000";
      s211 <= "0000000000000000000000000000000000";
      s212 <= "0000000000000000000000000000000000";
      s213 <= "0000000000000000000000000000000000";
      s214 <= "0000000000000000000000000000000000";
      s215 <= "0000000000000000000000000000000000";
      s216 <= "0000000000000000000000000000000000";
      s217 <= "0000000000000000000000000000000000";
      s218 <= "0000000000000000000000000000000000";
      s219 <= "0000000000000000000000000000000000";
      s220 <= "0000000000000000000000000000000000";
      s221 <= "0000000000000000000000000000000000";
      s222 <= "0000000000000000000000000000000000";
      s223 <= "0000000000000000000000000000000000";
      s224 <= "0000000000000000000000000000000000";
      s225 <= "0000000000000000000000000000000000";
      s226 <= "0000000000000000000000000000000000";
      s227 <= "0000000000000000000000000000000000";
      s228 <= "0000000000000000000000000000000000";
      s229 <= "0000000000000000000000000000000000";
      s230 <= "0000000000000000000000000000000000";
      s231 <= "0000000000000000000000000000000000";
      s232 <= "0000000000000000000000000000000000";
      s233 <= "0000000000000000000000000000000000";
      s234 <= "0000000000000000000000000000000000";
      s235 <= "0000000000000000000000000000000000";
      s236 <= "0000000000000000000000000000000000";
      s237 <= "0000000000000000000000000000000000";
      s238 <= "0000000000000000000000000000000000";
      s239 <= "0000000000000000000000000000000000";
      s240 <= "0000000000000000000000000000000000";
      s241 <= "0000000000000000000000000000000000";
      s242 <= "0000000000000000000000000000000000";
      s243 <= "0000000000000000000000000000000000";
      s244 <= "0000000000000000000000000000000000";
      s245 <= "0000000000000000000000000000000000";
      s246 <= "0000000000000000000000000000000000";
      s247 <= "0000000000000000000000000000000000";
      s248 <= "0000000000000000000000000000000000";
      s249 <= "0000000000000000000000000000000000";
      s250 <= "0000000000000000000000000000000000";
      s251 <= "0000000000000000000000000000000000";
      s252 <= "0000000000000000000000000000000000";
      s253 <= "0000000000000000000000000000000000";
      s254 <= "0000000000000000000000000000000000";
      s255 <= "0000000000000000000000000000000000";
      s256 <= "0000000000000000000000000000000000";
      s257 <= "0000000000000000000000000000000000";
      s258 <= "0000000000000000000000000000000000";
      s259 <= "0000000000000000000000000000000000";
      s260 <= "0000000000000000000000000000000000";
      s261 <= "0000000000000000000000000000000000";
      s262 <= "0000000000000000000000000000000000";
      s263 <= "0000000000000000000000000000000000";
      s264 <= "0000000000000000000000000000000000";
      s265 <= "0000000000000000000000000000000000";
      s266 <= "0000000000000000000000000000000000";
      s267 <= "0000000000000000000000000000000000";
      s268 <= "0000000000000000000000000000000000";
      s269 <= "0000000000000000000000000000000000";
      s270 <= "0000000000000000000000000000000000";
      s271 <= "0000000000000000000000000000000000";
      s272 <= "0000000000000000000000000000000000";
      s273 <= "0000000000000000000000000000000000";
      s274 <= "0000000000000000000000000000000000";
      s275 <= "0000000000000000000000000000000000";
      s276 <= "0000000000000000000000000000000000";
      s277 <= "0000000000000000000000000000000000";
      s278 <= "0000000000000000000000000000000000";
      s279 <= "0000000000000000000000000000000000";
      s280 <= "0000000000000000000000000000000000";
      s281 <= "0000000000000000000000000000000000";
      s282 <= "0000000000000000000000000000000000";
      s283 <= "0000000000000000000000000000000000";
      s284 <= "0000000000000000000000000000000000";
      s285 <= "0000000000000000000000000000000000";
      s286 <= "0000000000000000000000000000000000";
      s287 <= "0000000000000000000000000000000000";
      s288 <= "0000000000000000000000000000000000";
      s289 <= "0000000000000000000000000000000000";
      s290 <= "0000000000000000000000000000000000";
      s291 <= "0000000000000000000000000000000000";
      s292 <= "0000000000000000000000000000000000";
      s293 <= "0000000000000000000000000000000000";
      s294 <= "0000000000000000000000000000000000";
      s295 <= "0000000000000000000000000000000000";
      s296 <= "0000000000000000000000000000000000";
      s297 <= "0000000000000000000000000000000000";
      s298 <= "0000000000000000000000000000000000";
      s299 <= "0000000000000000000000000000000000";
      s300 <= "0000000000000000000000000000000000";
      s301 <= "0000000000000000000000000000000000";
      s302 <= "0000000000000000000000000000000000";
      s303 <= "0000000000000000000000000000000000";
      s304 <= "0000000000000000000000000000000000";
      s305 <= "0000000000000000000000000000000000";
      s306 <= "0000000000000000000000000000000000";
      s307 <= "0000000000000000000000000000000000";
      s308 <= "0000000000000000000000000000000000";
      s309 <= "0000000000000000000000000000000000";
      s310 <= "0000000000000000000000000000000000";
      s311 <= "0000000000000000000000000000000000";
      s312 <= "0000000000000000000000000000000000";
      s313 <= "0000000000000000000000000000000000";
      s314 <= "0000000000000000000000000000000000";
      s315 <= "0000000000000000000000000000000000";
      s316 <= "0000000000000000000000000000000000";
      s317 <= "0000000000000000000000000000000000";
      s318 <= "0000000000000000000000000000000000";
      s319 <= "0000000000000000000000000000000000";
      s320 <= "0000000000000000000000000000000000";
      s321 <= "0000000000000000000000000000000000";
      s322 <= "0000000000000000000000000000000000";
      s323 <= "0000000000000000000000000000000000";
      s324 <= "0000000000000000000000000000000000";
      s325 <= "0000000000000000000000000000000000";
      s326 <= "0000000000000000000000000000000000";
      s327 <= "0000000000000000000000000000000000";
      s328 <= "0000000000000000000000000000000000";
      s329 <= "0000000000000000000000000000000000";
      s330 <= "0000000000000000000000000000000000";
      s331 <= "0000000000000000000000000000000000";
      s332 <= "0000000000000000000000000000000000";
      s333 <= "0000000000000000000000000000000000";
      s334 <= "0000000000000000000000000000000000";
      s335 <= "0000000000000000000000000000000000";
      s336 <= "0000000000000000000000000000000000";
      s337 <= "0000000000000000000000000000000000";
      s338 <= "0000000000000000000000000000000000";
      s339 <= "0000000000000000000000000000000000";
      s340 <= "0000000000000000000000000000000000";
      s341 <= "0000000000000000000000000000000000";
      s342 <= "0000000000000000000000000000000000";
      s343 <= "0000000000000000000000000000000000";
      s344 <= "0000000000000000000000000000000000";
      s345 <= "0000000000000000000000000000000000";
      s346 <= "0000000000000000000000000000000000";
      s347 <= "0000000000000000000000000000000000";
      s348 <= "0000000000000000000000000000000000";
      s349 <= "0000000000000000000000000000000000";
      s350 <= "0000000000000000000000000000000000";
      s351 <= "0000000000000000000000000000000000";
      s352 <= "0000000000000000000000000000000000";
      s353 <= "0000000000000000000000000000000000";
      s354 <= "0000000000000000000000000000000000";
      s355 <= "0000000000000000000000000000000000";
      s356 <= "0000000000000000000000000000000000";
      s357 <= "0000000000000000000000000000000000";
      s358 <= "0000000000000000000000000000000000";
      s359 <= "0000000000000000000000000000000000";
      s360 <= "0000000000000000000000000000000000";
      s361 <= "0000000000000000000000000000000000";
      s362 <= "0000000000000000000000000000000000";
      s363 <= "0000000000000000000000000000000000";
      s364 <= "0000000000000000000000000000000000";
      s365 <= "0000000000000000000000000000000000";
      s366 <= "0000000000000000000000000000000000";
      s367 <= "0000000000000000000000000000000000";
      s368 <= "0000000000000000000000000000000000";
      s369 <= "0000000000000000000000000000000000";
      s370 <= "0000000000000000000000000000000000";
      s371 <= "0000000000000000000000000000000000";
      s372 <= "0000000000000000000000000000000000";
      s373 <= "0000000000000000000000000000000000";
      s374 <= "0000000000000000000000000000000000";
      s375 <= "0000000000000000000000000000000000";
      s376 <= "0000000000000000000000000000000000";
      s377 <= "0000000000000000000000000000000000";
      s378 <= "0000000000000000000000000000000000";
      s379 <= "0000000000000000000000000000000000";
      s380 <= "0000000000000000000000000000000000";
      s381 <= "0000000000000000000000000000000000";
      s382 <= "0000000000000000000000000000000000";
      s383 <= "0000000000000000000000000000000000";
      s384 <= "0000000000000000000000000000000000";
      s385 <= "0000000000000000000000000000000000";
      s386 <= "0000000000000000000000000000000000";
      s387 <= "0000000000000000000000000000000000";
      s388 <= "0000000000000000000000000000000000";
      s389 <= "0000000000000000000000000000000000";
      s390 <= "0000000000000000000000000000000000";
      s391 <= "0000000000000000000000000000000000";
      s392 <= "0000000000000000000000000000000000";
      s393 <= "0000000000000000000000000000000000";
      s394 <= "0000000000000000000000000000000000";
      s395 <= "0000000000000000000000000000000000";
      s396 <= "0000000000000000000000000000000000";
      s397 <= "0000000000000000000000000000000000";
      s398 <= "0000000000000000000000000000000000";
      s399 <= "0000000000000000000000000000000000";
      s400 <= "0000000000000000000000000000000000";
      s401 <= "0000000000000000000000000000000000";
      s402 <= "0000000000000000000000000000000000";
      s403 <= "0000000000000000000000000000000000";
      s404 <= "0000000000000000000000000000000000";
      s405 <= "0000000000000000000000000000000000";
      s406 <= "0000000000000000000000000000000000";
      s407 <= "0000000000000000000000000000000000";
      s408 <= "0000000000000000000000000000000000";
      s409 <= "0000000000000000000000000000000000";
      s410 <= "0000000000000000000000000000000000";
      s411 <= "0000000000000000000000000000000000";
      s412 <= "0000000000000000000000000000000000";
      s413 <= "0000000000000000000000000000000000";
      s414 <= "0000000000000000000000000000000000";
      s415 <= "0000000000000000000000000000000000";
      s416 <= "0000000000000000000000000000000000";
      s417 <= "0000000000000000000000000000000000";
      s418 <= "0000000000000000000000000000000000";
      s419 <= "0000000000000000000000000000000000";
      s420 <= "0000000000000000000000000000000000";
      s421 <= "0000000000000000000000000000000000";
      s422 <= "0000000000000000000000000000000000";
      s423 <= "0000000000000000000000000000000000";
      s424 <= "0000000000000000000000000000000000";
      s425 <= "0000000000000000000000000000000000";
      s426 <= "0000000000000000000000000000000000";
      s427 <= "0000000000000000000000000000000000";
      s428 <= "0000000000000000000000000000000000";
      s429 <= "0000000000000000000000000000000000";
      s430 <= "0000000000000000000000000000000000";
      s431 <= "0000000000000000000000000000000000";
      s432 <= "0000000000000000000000000000000000";
      s433 <= "0000000000000000000000000000000000";
      s434 <= "0000000000000000000000000000000000";
      s435 <= "0000000000000000000000000000000000";
      s436 <= "0000000000000000000000000000000000";
      s437 <= "0000000000000000000000000000000000";
      s438 <= "0000000000000000000000000000000000";
      s439 <= "0000000000000000000000000000000000";
      s440 <= "0000000000000000000000000000000000";
      s441 <= "0000000000000000000000000000000000";
      s442 <= "0000000000000000000000000000000000";
      s443 <= "0000000000000000000000000000000000";
      s444 <= "0000000000000000000000000000000000";
      s445 <= "0000000000000000000000000000000000";
      s446 <= "0000000000000000000000000000000000";
      s447 <= "0000000000000000000000000000000000";
      s448 <= "0000000000000000000000000000000000";
      s449 <= "0000000000000000000000000000000000";
      s450 <= "0000000000000000000000000000000000";
      s451 <= "0000000000000000000000000000000000";
      s452 <= "0000000000000000000000000000000000";
      s453 <= "0000000000000000000000000000000000";
      s454 <= "0000000000000000000000000000000000";
      s455 <= "0000000000000000000000000000000000";
      s456 <= "0000000000000000000000000000000000";
      s457 <= "0000000000000000000000000000000000";
      s458 <= "0000000000000000000000000000000000";
      s459 <= "0000000000000000000000000000000000";
      s460 <= "0000000000000000000000000000000000";
      s461 <= "0000000000000000000000000000000000";
      s462 <= "0000000000000000000000000000000000";
      s463 <= "0000000000000000000000000000000000";
      s464 <= "0000000000000000000000000000000000";
      s465 <= "0000000000000000000000000000000000";
      s466 <= "0000000000000000000000000000000000";
      s467 <= "0000000000000000000000000000000000";
      s468 <= "0000000000000000000000000000000000";
      s469 <= "0000000000000000000000000000000000";
      s470 <= "0000000000000000000000000000000000";
      s471 <= "0000000000000000000000000000000000";
      s472 <= "0000000000000000000000000000000000";
      s473 <= "0000000000000000000000000000000000";
      s474 <= "0000000000000000000000000000000000";
      s475 <= "0000000000000000000000000000000000";
      s476 <= "0000000000000000000000000000000000";
      s477 <= "0000000000000000000000000000000000";
      s478 <= "0000000000000000000000000000000000";
      s479 <= "0000000000000000000000000000000000";
      s480 <= "0000000000000000000000000000000000";
      s481 <= "0000000000000000000000000000000000";
      s482 <= "0000000000000000000000000000000000";
      s483 <= "0000000000000000000000000000000000";
      s484 <= "0000000000000000000000000000000000";
      s485 <= "0000000000000000000000000000000000";
      s486 <= "0000000000000000000000000000000000";
      s487 <= "0000000000000000000000000000000000";
      s488 <= "0000000000000000000000000000000000";
      s489 <= "0000000000000000000000000000000000";
      s490 <= "0000000000000000000000000000000000";
      s491 <= "0000000000000000000000000000000000";
      s492 <= "0000000000000000000000000000000000";
      s493 <= "0000000000000000000000000000000000";
      s494 <= "0000000000000000000000000000000000";
      s495 <= "0000000000000000000000000000000000";
      s496 <= "0000000000000000000000000000000000";
      s497 <= "0000000000000000000000000000000000";
      s498 <= "0000000000000000000000000000000000";
      s499 <= "0000000000000000000000000000000000";
      s500 <= "0000000000000000000000000000000000";
      s501 <= "0000000000000000000000000000000000";
      s502 <= "0000000000000000000000000000000000";
      s503 <= "0000000000000000000000000000000000";
      s504 <= "0000000000000000000000000000000000";
      s505 <= "0000000000000000000000000000000000";
      s506 <= "0000000000000000000000000000000000";
      s507 <= "0000000000000000000000000000000000";
      s508 <= "0000000000000000000000000000000000";
      s509 <= "0000000000000000000000000000000000";
      s510 <= "0000000000000000000000000000000000";
      s511 <= "0000000000000000000000000000000000";
      s512 <= "0000000000000000000000000000000000";
      s513 <= "0000000000000000000000000000000000";
      s514 <= "0000000000000000000000000000000000";
      s515 <= "0000000000000000000000000000000000";
      s516 <= "0000000000000000000000000000000000";
      s517 <= "0000000000000000000000000000000000";
      s518 <= "0000000000000000000000000000000000";
      s519 <= "0000000000000000000000000000000000";
      s520 <= "0000000000000000000000000000000000";
      s521 <= "0000000000000000000000000000000000";
      s522 <= "0000000000000000000000000000000000";
      s523 <= "0000000000000000000000000000000000";
      s524 <= "0000000000000000000000000000000000";
      s525 <= "0000000000000000000000000000000000";
      s526 <= "0000000000000000000000000000000000";
      s527 <= "0000000000000000000000000000000000";
      s528 <= "0000000000000000000000000000000000";
      s529 <= "0000000000000000000000000000000000";
      s530 <= "0000000000000000000000000000000000";
      s531 <= "0000000000000000000000000000000000";
      s532 <= "0000000000000000000000000000000000";
      s533 <= "0000000000000000000000000000000000";
      s534 <= "0000000000000000000000000000000000";
      s535 <= "0000000000000000000000000000000000";
      s536 <= "0000000000000000000000000000000000";
      s537 <= "0000000000000000000000000000000000";
      s538 <= "0000000000000000000000000000000000";
      s539 <= "0000000000000000000000000000000000";
      s540 <= "0000000000000000000000000000000000";
      s541 <= "0000000000000000000000000000000000";
      s542 <= "0000000000000000000000000000000000";
      s543 <= "0000000000000000000000000000000000";
      s544 <= "0000000000000000000000000000000000";
      s545 <= "0000000000000000000000000000000000";
      s546 <= "0000000000000000000000000000000000";
      s547 <= "0000000000000000000000000000000000";
      s548 <= "0000000000000000000000000000000000";
      s549 <= "0000000000000000000000000000000000";
      s550 <= "0000000000000000000000000000000000";
      s551 <= "0000000000000000000000000000000000";
      s552 <= "0000000000000000000000000000000000";
      s553 <= "0000000000000000000000000000000000";
      s554 <= "0000000000000000000000000000000000";
      s555 <= "0000000000000000000000000000000000";
      s556 <= "0000000000000000000000000000000000";
      s557 <= "0000000000000000000000000000000000";
      s558 <= "0000000000000000000000000000000000";
      s559 <= "0000000000000000000000000000000000";
      s560 <= "0000000000000000000000000000000000";
      s561 <= "0000000000000000000000000000000000";
      s562 <= "0000000000000000000000000000000000";
      s563 <= "0000000000000000000000000000000000";
      s564 <= "0000000000000000000000000000000000";
      s565 <= "0000000000000000000000000000000000";
      s566 <= "0000000000000000000000000000000000";
      s567 <= "0000000000000000000000000000000000";
      s568 <= "0000000000000000000000000000000000";
      s569 <= "0000000000000000000000000000000000";
      s570 <= "0000000000000000000000000000000000";
      s571 <= "0000000000000000000000000000000000";
      s572 <= "0000000000000000000000000000000000";
      s573 <= "0000000000000000000000000000000000";
      s574 <= "0000000000000000000000000000000000";
      s575 <= "0000000000000000000000000000000000";
      s576 <= "0000000000000000000000000000000000";
      s577 <= "0000000000000000000000000000000000";
      s578 <= "0000000000000000000000000000000000";
      s579 <= "0000000000000000000000000000000000";
      s580 <= "0000000000000000000000000000000000";
      s581 <= "0000000000000000000000000000000000";
      s582 <= "0000000000000000000000000000000000";
      s583 <= "0000000000000000000000000000000000";
      s584 <= "0000000000000000000000000000000000";
      s585 <= "0000000000000000000000000000000000";
      s586 <= "0000000000000000000000000000000000";
      s587 <= "0000000000000000000000000000000000";
      s588 <= "0000000000000000000000000000000000";
      s589 <= "0000000000000000000000000000000000";
      s590 <= "0000000000000000000000000000000000";
      s591 <= "0000000000000000000000000000000000";
      s592 <= "0000000000000000000000000000000000";
      s593 <= "0000000000000000000000000000000000";
      s594 <= "0000000000000000000000000000000000";
      s595 <= "0000000000000000000000000000000000";
      s596 <= "0000000000000000000000000000000000";
      s597 <= "0000000000000000000000000000000000";
      s598 <= "0000000000000000000000000000000000";
      s599 <= "0000000000000000000000000000000000";
      s600 <= "0000000000000000000000000000000000";
      s601 <= "0000000000000000000000000000000000";
      s602 <= "0000000000000000000000000000000000";
      s603 <= "0000000000000000000000000000000000";
      s604 <= "0000000000000000000000000000000000";
      s605 <= "0000000000000000000000000000000000";
      s606 <= "0000000000000000000000000000000000";
      s607 <= "0000000000000000000000000000000000";
      s608 <= "0000000000000000000000000000000000";
      s609 <= "0000000000000000000000000000000000";
      s610 <= "0000000000000000000000000000000000";
      s611 <= "0000000000000000000000000000000000";
      s612 <= "0000000000000000000000000000000000";
      s613 <= "0000000000000000000000000000000000";
      s614 <= "0000000000000000000000000000000000";
      s615 <= "0000000000000000000000000000000000";
      s616 <= "0000000000000000000000000000000000";
      s617 <= "0000000000000000000000000000000000";
      s618 <= "0000000000000000000000000000000000";
      s619 <= "0000000000000000000000000000000000";
      s620 <= "0000000000000000000000000000000000";
      s621 <= "0000000000000000000000000000000000";
      s622 <= "0000000000000000000000000000000000";
      s623 <= "0000000000000000000000000000000000";
      s624 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      s165 <= s164;
      s166 <= s165;
      s167 <= s166;
      s168 <= s167;
      s169 <= s168;
      s170 <= s169;
      s171 <= s170;
      s172 <= s171;
      s173 <= s172;
      s174 <= s173;
      s175 <= s174;
      s176 <= s175;
      s177 <= s176;
      s178 <= s177;
      s179 <= s178;
      s180 <= s179;
      s181 <= s180;
      s182 <= s181;
      s183 <= s182;
      s184 <= s183;
      s185 <= s184;
      s186 <= s185;
      s187 <= s186;
      s188 <= s187;
      s189 <= s188;
      s190 <= s189;
      s191 <= s190;
      s192 <= s191;
      s193 <= s192;
      s194 <= s193;
      s195 <= s194;
      s196 <= s195;
      s197 <= s196;
      s198 <= s197;
      s199 <= s198;
      s200 <= s199;
      s201 <= s200;
      s202 <= s201;
      s203 <= s202;
      s204 <= s203;
      s205 <= s204;
      s206 <= s205;
      s207 <= s206;
      s208 <= s207;
      s209 <= s208;
      s210 <= s209;
      s211 <= s210;
      s212 <= s211;
      s213 <= s212;
      s214 <= s213;
      s215 <= s214;
      s216 <= s215;
      s217 <= s216;
      s218 <= s217;
      s219 <= s218;
      s220 <= s219;
      s221 <= s220;
      s222 <= s221;
      s223 <= s222;
      s224 <= s223;
      s225 <= s224;
      s226 <= s225;
      s227 <= s226;
      s228 <= s227;
      s229 <= s228;
      s230 <= s229;
      s231 <= s230;
      s232 <= s231;
      s233 <= s232;
      s234 <= s233;
      s235 <= s234;
      s236 <= s235;
      s237 <= s236;
      s238 <= s237;
      s239 <= s238;
      s240 <= s239;
      s241 <= s240;
      s242 <= s241;
      s243 <= s242;
      s244 <= s243;
      s245 <= s244;
      s246 <= s245;
      s247 <= s246;
      s248 <= s247;
      s249 <= s248;
      s250 <= s249;
      s251 <= s250;
      s252 <= s251;
      s253 <= s252;
      s254 <= s253;
      s255 <= s254;
      s256 <= s255;
      s257 <= s256;
      s258 <= s257;
      s259 <= s258;
      s260 <= s259;
      s261 <= s260;
      s262 <= s261;
      s263 <= s262;
      s264 <= s263;
      s265 <= s264;
      s266 <= s265;
      s267 <= s266;
      s268 <= s267;
      s269 <= s268;
      s270 <= s269;
      s271 <= s270;
      s272 <= s271;
      s273 <= s272;
      s274 <= s273;
      s275 <= s274;
      s276 <= s275;
      s277 <= s276;
      s278 <= s277;
      s279 <= s278;
      s280 <= s279;
      s281 <= s280;
      s282 <= s281;
      s283 <= s282;
      s284 <= s283;
      s285 <= s284;
      s286 <= s285;
      s287 <= s286;
      s288 <= s287;
      s289 <= s288;
      s290 <= s289;
      s291 <= s290;
      s292 <= s291;
      s293 <= s292;
      s294 <= s293;
      s295 <= s294;
      s296 <= s295;
      s297 <= s296;
      s298 <= s297;
      s299 <= s298;
      s300 <= s299;
      s301 <= s300;
      s302 <= s301;
      s303 <= s302;
      s304 <= s303;
      s305 <= s304;
      s306 <= s305;
      s307 <= s306;
      s308 <= s307;
      s309 <= s308;
      s310 <= s309;
      s311 <= s310;
      s312 <= s311;
      s313 <= s312;
      s314 <= s313;
      s315 <= s314;
      s316 <= s315;
      s317 <= s316;
      s318 <= s317;
      s319 <= s318;
      s320 <= s319;
      s321 <= s320;
      s322 <= s321;
      s323 <= s322;
      s324 <= s323;
      s325 <= s324;
      s326 <= s325;
      s327 <= s326;
      s328 <= s327;
      s329 <= s328;
      s330 <= s329;
      s331 <= s330;
      s332 <= s331;
      s333 <= s332;
      s334 <= s333;
      s335 <= s334;
      s336 <= s335;
      s337 <= s336;
      s338 <= s337;
      s339 <= s338;
      s340 <= s339;
      s341 <= s340;
      s342 <= s341;
      s343 <= s342;
      s344 <= s343;
      s345 <= s344;
      s346 <= s345;
      s347 <= s346;
      s348 <= s347;
      s349 <= s348;
      s350 <= s349;
      s351 <= s350;
      s352 <= s351;
      s353 <= s352;
      s354 <= s353;
      s355 <= s354;
      s356 <= s355;
      s357 <= s356;
      s358 <= s357;
      s359 <= s358;
      s360 <= s359;
      s361 <= s360;
      s362 <= s361;
      s363 <= s362;
      s364 <= s363;
      s365 <= s364;
      s366 <= s365;
      s367 <= s366;
      s368 <= s367;
      s369 <= s368;
      s370 <= s369;
      s371 <= s370;
      s372 <= s371;
      s373 <= s372;
      s374 <= s373;
      s375 <= s374;
      s376 <= s375;
      s377 <= s376;
      s378 <= s377;
      s379 <= s378;
      s380 <= s379;
      s381 <= s380;
      s382 <= s381;
      s383 <= s382;
      s384 <= s383;
      s385 <= s384;
      s386 <= s385;
      s387 <= s386;
      s388 <= s387;
      s389 <= s388;
      s390 <= s389;
      s391 <= s390;
      s392 <= s391;
      s393 <= s392;
      s394 <= s393;
      s395 <= s394;
      s396 <= s395;
      s397 <= s396;
      s398 <= s397;
      s399 <= s398;
      s400 <= s399;
      s401 <= s400;
      s402 <= s401;
      s403 <= s402;
      s404 <= s403;
      s405 <= s404;
      s406 <= s405;
      s407 <= s406;
      s408 <= s407;
      s409 <= s408;
      s410 <= s409;
      s411 <= s410;
      s412 <= s411;
      s413 <= s412;
      s414 <= s413;
      s415 <= s414;
      s416 <= s415;
      s417 <= s416;
      s418 <= s417;
      s419 <= s418;
      s420 <= s419;
      s421 <= s420;
      s422 <= s421;
      s423 <= s422;
      s424 <= s423;
      s425 <= s424;
      s426 <= s425;
      s427 <= s426;
      s428 <= s427;
      s429 <= s428;
      s430 <= s429;
      s431 <= s430;
      s432 <= s431;
      s433 <= s432;
      s434 <= s433;
      s435 <= s434;
      s436 <= s435;
      s437 <= s436;
      s438 <= s437;
      s439 <= s438;
      s440 <= s439;
      s441 <= s440;
      s442 <= s441;
      s443 <= s442;
      s444 <= s443;
      s445 <= s444;
      s446 <= s445;
      s447 <= s446;
      s448 <= s447;
      s449 <= s448;
      s450 <= s449;
      s451 <= s450;
      s452 <= s451;
      s453 <= s452;
      s454 <= s453;
      s455 <= s454;
      s456 <= s455;
      s457 <= s456;
      s458 <= s457;
      s459 <= s458;
      s460 <= s459;
      s461 <= s460;
      s462 <= s461;
      s463 <= s462;
      s464 <= s463;
      s465 <= s464;
      s466 <= s465;
      s467 <= s466;
      s468 <= s467;
      s469 <= s468;
      s470 <= s469;
      s471 <= s470;
      s472 <= s471;
      s473 <= s472;
      s474 <= s473;
      s475 <= s474;
      s476 <= s475;
      s477 <= s476;
      s478 <= s477;
      s479 <= s478;
      s480 <= s479;
      s481 <= s480;
      s482 <= s481;
      s483 <= s482;
      s484 <= s483;
      s485 <= s484;
      s486 <= s485;
      s487 <= s486;
      s488 <= s487;
      s489 <= s488;
      s490 <= s489;
      s491 <= s490;
      s492 <= s491;
      s493 <= s492;
      s494 <= s493;
      s495 <= s494;
      s496 <= s495;
      s497 <= s496;
      s498 <= s497;
      s499 <= s498;
      s500 <= s499;
      s501 <= s500;
      s502 <= s501;
      s503 <= s502;
      s504 <= s503;
      s505 <= s504;
      s506 <= s505;
      s507 <= s506;
      s508 <= s507;
      s509 <= s508;
      s510 <= s509;
      s511 <= s510;
      s512 <= s511;
      s513 <= s512;
      s514 <= s513;
      s515 <= s514;
      s516 <= s515;
      s517 <= s516;
      s518 <= s517;
      s519 <= s518;
      s520 <= s519;
      s521 <= s520;
      s522 <= s521;
      s523 <= s522;
      s524 <= s523;
      s525 <= s524;
      s526 <= s525;
      s527 <= s526;
      s528 <= s527;
      s529 <= s528;
      s530 <= s529;
      s531 <= s530;
      s532 <= s531;
      s533 <= s532;
      s534 <= s533;
      s535 <= s534;
      s536 <= s535;
      s537 <= s536;
      s538 <= s537;
      s539 <= s538;
      s540 <= s539;
      s541 <= s540;
      s542 <= s541;
      s543 <= s542;
      s544 <= s543;
      s545 <= s544;
      s546 <= s545;
      s547 <= s546;
      s548 <= s547;
      s549 <= s548;
      s550 <= s549;
      s551 <= s550;
      s552 <= s551;
      s553 <= s552;
      s554 <= s553;
      s555 <= s554;
      s556 <= s555;
      s557 <= s556;
      s558 <= s557;
      s559 <= s558;
      s560 <= s559;
      s561 <= s560;
      s562 <= s561;
      s563 <= s562;
      s564 <= s563;
      s565 <= s564;
      s566 <= s565;
      s567 <= s566;
      s568 <= s567;
      s569 <= s568;
      s570 <= s569;
      s571 <= s570;
      s572 <= s571;
      s573 <= s572;
      s574 <= s573;
      s575 <= s574;
      s576 <= s575;
      s577 <= s576;
      s578 <= s577;
      s579 <= s578;
      s580 <= s579;
      s581 <= s580;
      s582 <= s581;
      s583 <= s582;
      s584 <= s583;
      s585 <= s584;
      s586 <= s585;
      s587 <= s586;
      s588 <= s587;
      s589 <= s588;
      s590 <= s589;
      s591 <= s590;
      s592 <= s591;
      s593 <= s592;
      s594 <= s593;
      s595 <= s594;
      s596 <= s595;
      s597 <= s596;
      s598 <= s597;
      s599 <= s598;
      s600 <= s599;
      s601 <= s600;
      s602 <= s601;
      s603 <= s602;
      s604 <= s603;
      s605 <= s604;
      s606 <= s605;
      s607 <= s606;
      s608 <= s607;
      s609 <= s608;
      s610 <= s609;
      s611 <= s610;
      s612 <= s611;
      s613 <= s612;
      s614 <= s613;
      s615 <= s614;
      s616 <= s615;
      s617 <= s616;
      s618 <= s617;
      s619 <= s618;
      s620 <= s619;
      s621 <= s620;
      s622 <= s621;
      s623 <= s622;
      s624 <= s623;
      Y <= s624;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 60 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      Y <= s59;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 69 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      Y <= s68;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          In2_0 : in std_logic_vector(31 downto 0);
          Out2_0 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_64_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(5 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_64_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iS_51 : in std_logic_vector(33 downto 0);
             iS_52 : in std_logic_vector(33 downto 0);
             iS_53 : in std_logic_vector(33 downto 0);
             iS_54 : in std_logic_vector(33 downto 0);
             iS_55 : in std_logic_vector(33 downto 0);
             iS_56 : in std_logic_vector(33 downto 0);
             iS_57 : in std_logic_vector(33 downto 0);
             iS_58 : in std_logic_vector(33 downto 0);
             iS_59 : in std_logic_vector(33 downto 0);
             iS_60 : in std_logic_vector(33 downto 0);
             iS_61 : in std_logic_vector(33 downto 0);
             iS_62 : in std_logic_vector(33 downto 0);
             iS_63 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_61_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iS_51 : in std_logic_vector(33 downto 0);
             iS_52 : in std_logic_vector(33 downto 0);
             iS_53 : in std_logic_vector(33 downto 0);
             iS_54 : in std_logic_vector(33 downto 0);
             iS_55 : in std_logic_vector(33 downto 0);
             iS_56 : in std_logic_vector(33 downto 0);
             iS_57 : in std_logic_vector(33 downto 0);
             iS_58 : in std_logic_vector(33 downto 0);
             iS_59 : in std_logic_vector(33 downto 0);
             iS_60 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_34_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_51_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_20_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(4 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_13_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_6_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_3_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(1 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_2_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(0 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_0_617123672897668340553423149685841053724_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_631862801488796588245122620719484984875_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_436934552725145586293820088030770421028_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_561088850170149200380365073215216398239_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_67381401040949318037576176720904186368_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_767419732788928943278961014584638178349_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_83466961525726479642628419242100790143_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_869869533302351394254969818575773388147_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_663686724095854829741369940165895968676_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_712333225863809871292176012502750381827_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_777424256340159325340266605053329840302_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_858338451424324633265428019512910395861_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_95403875322976861017565397560247220099_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_062858000783881262663044253713451325893_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_182256984960216694702239692560397088528_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_308589307952890523623068474989850074053_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_99584180311675085661704542872030287981_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_987534845729581944873132215434452518821_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_906979034015293006376623452524654567242_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_898568629504465254953515795932617038488_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_891139475905879052675118145998567342758_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_885091234632599865861379839770961552858_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_880803415623673480183697392931208014488_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_878576235602384070233483726042322814465_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_979173278459382512295405831537209451199_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_970685163049390786760284299816703423858_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_962013487567665803723571116279345005751_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_95312319664069156122110371143207885325_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_944010225685960935315677033941028639674_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_934712586109242460352675152535084635019_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_925322845902050161726037913467735052109_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n0_916000226493365876656582713621901348233_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum1_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum1_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum1_1_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum1_1_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum1_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum1_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum12_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum12_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum15_2_impl_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum15_2_impl_1_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum2_2_impl_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum2_2_impl_1_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum26_1_impl_0_LUT_wIn_6_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum26_1_impl_1_LUT_wIn_6_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum41_2_impl_0_LUT_wIn_6_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum41_2_impl_1_LUT_wIn_6_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum42_2_impl_0_LUT_wIn_6_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Sum42_2_impl_1_LUT_wIn_6_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Out2_0_0_LUT_wIn_6_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_100_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_684_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_746_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_849_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_948_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1016_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1081_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_162_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_246_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_296_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_365_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_439_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_507_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_558_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_624_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_73_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_75_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_70_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_130_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_681_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_735_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_838_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_946_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_995_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1056_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_146_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_239_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_294_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_359_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_442_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_499_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_555_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_625_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount641_out : std_logic_vector(5 downto 0) := (others => '0');
signal In2_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum1_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum1_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum1_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum1_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum1_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum1_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum1_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum1_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum15_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum15_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum15_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum26_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum26_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum26_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum41_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum41_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum41_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum42_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum42_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum42_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal a_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a10_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a14_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a15_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a3_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a8_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal a9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal b_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c10_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c14_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c15_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c3_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c8_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal c9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal d_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Out2_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay57No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay60No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay63No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay63No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay62No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay71No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay67No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay66No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum1_0_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Sum1_0_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Sum1_1_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Sum1_1_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Sum1_2_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Sum1_2_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Sum12_2_impl_0_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Sum12_2_impl_1_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Sum15_2_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Sum15_2_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Sum2_2_impl_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Sum2_2_impl_1_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Sum26_1_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Sum26_1_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Sum41_2_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Sum41_2_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Sum42_2_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Sum42_2_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Out2_0_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal In2_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No_out_to_Product_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out_to_Product_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay67No1_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay71No1_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay63No3_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out_to_Product_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out_to_Product_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay66No2_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay60No_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay62No4_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out_to_Product_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out_to_Product_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay63No2_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out_to_Sum1_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out_to_Sum1_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay57No2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out_to_Sum1_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out_to_Sum1_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out_to_Sum1_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out_to_Sum1_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No2_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out_to_Sum12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out_to_Sum12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out_to_Sum15_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out_to_Sum15_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out_to_Sum2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out_to_Sum2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out_to_Sum26_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out_to_Sum26_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Sum26_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Sum26_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Sum26_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Sum26_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum26_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Sum26_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out_to_Sum41_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out_to_Sum41_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Sum41_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Sum41_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Sum41_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Sum41_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out_to_Sum42_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out_to_Sum42_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Sum42_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Sum42_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Sum42_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Sum42_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Out2_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Out2_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Out2_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Out2_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount641_instance: ModuloCounter_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount641_out);
In2_0_IEEE <= In2_0;
   In2_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => In2_0_out,
                 X => In2_0_IEEE);

Delay1No_out_to_Product_0_impl_parent_implementedSystem_port_0_cast <= Delay1No_out;
Delay1No1_out_to_Product_0_impl_parent_implementedSystem_port_1_cast <= Delay1No1_out;
   Product_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product_0_impl_out,
                 X => Delay1No_out_to_Product_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No1_out_to_Product_0_impl_parent_implementedSystem_port_1_cast);

SharedReg271_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg271_out;
SharedReg304_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg304_out;
SharedReg273_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg273_out;
SharedReg305_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg305_out;
SharedReg274_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg274_out;
SharedReg306_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg306_out;
SharedReg289_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg289_out;
SharedReg307_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg307_out;
SharedReg308_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg308_out;
SharedReg269_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg269_out;
SharedReg275_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg275_out;
SharedReg272_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg272_out;
SharedReg276_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg276_out;
SharedReg277_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg277_out;
SharedReg309_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg309_out;
SharedReg310_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg310_out;
SharedReg278_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg278_out;
SharedReg257_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg257_out;
SharedReg293_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg293_out;
SharedReg279_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg279_out;
SharedReg311_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg311_out;
SharedReg280_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg280_out;
SharedReg312_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg312_out;
SharedReg281_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg281_out;
SharedReg313_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg313_out;
SharedReg282_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg282_out;
SharedReg314_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg314_out;
SharedReg283_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg283_out;
SharedReg315_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg315_out;
SharedReg284_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg284_out;
SharedReg316_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg316_out;
SharedReg288_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg288_out;
SharedReg292_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg292_out;
SharedReg286_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg286_out;
SharedReg261_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg261_out;
SharedReg291_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg291_out;
SharedReg254_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg254_out;
SharedReg285_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg285_out;
SharedReg295_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg295_out;
SharedReg296_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg296_out;
SharedReg263_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg263_out;
SharedReg287_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg287_out;
SharedReg256_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg256_out;
SharedReg299_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg299_out;
SharedReg255_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg255_out;
SharedReg264_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg264_out;
SharedReg267_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg267_out;
SharedReg294_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg294_out;
SharedReg268_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg268_out;
SharedReg300_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg300_out;
SharedReg290_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg290_out;
SharedReg298_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg298_out;
SharedReg258_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg258_out;
SharedReg253_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg253_out;
SharedReg262_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg262_out;
SharedReg265_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg265_out;
SharedReg259_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg259_out;
SharedReg260_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg260_out;
SharedReg297_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg297_out;
SharedReg266_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_60_cast <= SharedReg266_out;
SharedReg301_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_61_cast <= SharedReg301_out;
SharedReg302_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_62_cast <= SharedReg302_out;
SharedReg270_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_63_cast <= SharedReg270_out;
SharedReg303_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_64_cast <= SharedReg303_out;
   MUX_Product_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg271_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg304_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg275_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg272_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg276_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg277_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg309_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg310_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg278_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg257_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg293_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg279_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg273_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg311_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg280_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg312_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg281_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg313_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg282_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg314_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg283_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg315_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg284_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg305_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg316_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg288_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg292_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg286_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg261_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg291_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg254_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg285_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg295_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg296_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg274_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg263_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg287_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg256_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg299_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg255_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg264_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg267_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg294_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg268_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg300_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg306_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg290_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg298_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg258_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg253_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg262_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg265_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg259_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg260_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg297_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg266_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg289_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg301_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg302_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg270_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg303_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg307_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg308_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg269_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product_0_impl_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_0_impl_0_out,
                 Y => Delay1No_out);

SharedReg154_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg154_out;
SharedReg157_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg157_out;
SharedReg118_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg118_out;
SharedReg196_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg196_out;
SharedReg188_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg188_out;
SharedReg90_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg90_out;
SharedReg65_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg65_out;
SharedReg123_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg123_out;
SharedReg213_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg213_out;
SharedReg226_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg226_out;
SharedReg205_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg205_out;
SharedReg73_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg73_out;
SharedReg241_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg241_out;
SharedReg231_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg231_out;
SharedReg129_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg129_out;
SharedReg170_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg170_out;
SharedReg84_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg84_out;
SharedReg197_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg197_out;
SharedReg106_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg106_out;
SharedReg211_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg211_out;
SharedReg172_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg172_out;
SharedReg124_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg124_out;
Delay67No1_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_23_cast <= Delay67No1_out;
Delay71No1_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_24_cast <= Delay71No1_out;
SharedReg81_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg81_out;
SharedReg248_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg248_out;
SharedReg235_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg235_out;
SharedReg252_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg252_out;
Delay63No3_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_29_cast <= Delay63No3_out;
SharedReg164_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg164_out;
SharedReg174_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg174_out;
SharedReg141_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg141_out;
SharedReg134_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg134_out;
SharedReg112_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg112_out;
SharedReg131_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg131_out;
SharedReg237_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg237_out;
SharedReg131_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg131_out;
SharedReg180_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg180_out;
SharedReg188_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg188_out;
SharedReg69_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg69_out;
SharedReg104_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg104_out;
SharedReg145_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg145_out;
SharedReg100_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg100_out;
SharedReg113_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg113_out;
SharedReg197_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg197_out;
SharedReg176_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg176_out;
SharedReg220_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg220_out;
SharedReg143_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg143_out;
SharedReg58_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg58_out;
SharedReg148_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg148_out;
SharedReg225_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg225_out;
SharedReg204_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg204_out;
SharedReg245_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg245_out;
SharedReg219_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg219_out;
SharedReg58_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg58_out;
SharedReg198_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg198_out;
SharedReg249_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg249_out;
SharedReg137_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg137_out;
SharedReg117_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg117_out;
SharedReg238_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_60_cast <= SharedReg238_out;
SharedReg189_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_61_cast <= SharedReg189_out;
SharedReg125_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_62_cast <= SharedReg125_out;
SharedReg151_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_63_cast <= SharedReg151_out;
SharedReg127_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_64_cast <= SharedReg127_out;
   MUX_Product_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg154_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg157_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg205_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg73_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg241_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg231_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg129_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg170_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg84_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg197_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg106_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg211_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg118_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg172_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg124_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => Delay67No1_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => Delay71No1_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg81_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg248_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg235_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg252_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => Delay63No3_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg164_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg196_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg174_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg141_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg134_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg112_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg131_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg237_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg131_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg180_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg188_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg69_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg188_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg104_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg145_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg100_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg113_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg197_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg176_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg220_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg143_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg58_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg148_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg90_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg225_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg204_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg245_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg219_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg58_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg198_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg249_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg137_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg117_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg238_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg65_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg189_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg125_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg151_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg127_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg123_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg213_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg226_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product_0_impl_1_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_0_impl_1_out,
                 Y => Delay1No1_out);

Delay1No2_out_to_Product_1_impl_parent_implementedSystem_port_0_cast <= Delay1No2_out;
Delay1No3_out_to_Product_1_impl_parent_implementedSystem_port_1_cast <= Delay1No3_out;
   Product_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product_1_impl_out,
                 X => Delay1No2_out_to_Product_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No3_out_to_Product_1_impl_parent_implementedSystem_port_1_cast);

SharedReg299_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg299_out;
SharedReg255_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg255_out;
SharedReg264_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg264_out;
SharedReg267_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg267_out;
SharedReg294_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg294_out;
SharedReg268_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg268_out;
SharedReg300_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg300_out;
SharedReg290_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg290_out;
SharedReg298_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg298_out;
SharedReg258_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg258_out;
SharedReg253_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg253_out;
SharedReg262_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg262_out;
SharedReg265_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg265_out;
SharedReg259_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg259_out;
SharedReg260_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg260_out;
SharedReg297_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg297_out;
SharedReg266_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg266_out;
SharedReg301_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg301_out;
SharedReg302_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg302_out;
SharedReg270_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg270_out;
SharedReg303_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg303_out;
SharedReg271_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg271_out;
SharedReg304_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg304_out;
SharedReg273_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg273_out;
SharedReg305_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg305_out;
SharedReg274_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg274_out;
SharedReg306_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg306_out;
SharedReg289_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg289_out;
SharedReg307_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg307_out;
SharedReg308_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg308_out;
SharedReg269_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg269_out;
SharedReg275_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg275_out;
SharedReg272_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg272_out;
SharedReg276_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg276_out;
SharedReg277_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg277_out;
SharedReg309_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg309_out;
SharedReg310_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg310_out;
SharedReg278_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg278_out;
SharedReg257_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg257_out;
SharedReg293_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg293_out;
SharedReg279_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg279_out;
SharedReg311_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg311_out;
SharedReg280_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg280_out;
SharedReg312_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg312_out;
SharedReg281_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg281_out;
SharedReg313_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg313_out;
SharedReg282_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg282_out;
SharedReg314_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg314_out;
SharedReg283_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg283_out;
SharedReg315_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg315_out;
SharedReg284_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg284_out;
SharedReg316_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg316_out;
SharedReg288_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg288_out;
SharedReg292_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg292_out;
SharedReg286_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg286_out;
SharedReg261_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg261_out;
SharedReg291_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg291_out;
SharedReg254_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg254_out;
SharedReg285_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg285_out;
SharedReg295_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg295_out;
SharedReg296_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg296_out;
SharedReg263_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg263_out;
SharedReg287_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg287_out;
SharedReg256_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg256_out;
   MUX_Product_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg299_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg255_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg253_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg262_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg265_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg259_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg260_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg297_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg266_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg301_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg302_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg270_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg264_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg303_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg271_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg304_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg273_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg305_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg274_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg306_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg289_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg307_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg308_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg267_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg269_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg275_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg272_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg276_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg277_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg309_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg310_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg278_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg257_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg293_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg294_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg279_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg311_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg280_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg312_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg281_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg313_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg282_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg314_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg283_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg315_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg268_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg284_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg316_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg288_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg292_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg286_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg261_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg291_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg254_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg285_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg295_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg300_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg296_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg263_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg287_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg256_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg290_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg298_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg258_out_to_MUX_Product_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product_1_impl_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_1_impl_0_out,
                 Y => Delay1No2_out);

SharedReg225_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg225_out;
SharedReg131_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg131_out;
SharedReg59_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg59_out;
SharedReg102_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg102_out;
SharedReg67_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg67_out;
SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg58_out;
SharedReg74_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg74_out;
SharedReg246_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg246_out;
SharedReg240_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg240_out;
SharedReg197_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg197_out;
SharedReg101_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg101_out;
SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg58_out;
SharedReg134_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg134_out;
SharedReg221_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg221_out;
SharedReg63_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg63_out;
SharedReg208_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg208_out;
SharedReg180_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg180_out;
SharedReg230_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg230_out;
SharedReg167_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg167_out;
SharedReg78_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg78_out;
SharedReg169_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg169_out;
SharedReg82_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg82_out;
SharedReg84_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg84_out;
SharedReg154_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg154_out;
SharedReg128_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg128_out;
SharedReg76_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg76_out;
SharedReg195_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg195_out;
SharedReg200_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg200_out;
SharedReg212_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg212_out;
SharedReg244_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg244_out;
SharedReg113_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg113_out;
SharedReg147_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg147_out;
SharedReg73_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg73_out;
SharedReg188_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg188_out;
SharedReg121_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg121_out;
SharedReg234_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg234_out;
SharedReg92_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg92_out;
SharedReg84_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg84_out;
SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg58_out;
SharedReg136_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg136_out;
SharedReg161_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg161_out;
SharedReg217_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg217_out;
SharedReg88_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg88_out;
Delay66No2_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_44_cast <= Delay66No2_out;
SharedReg99_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg99_out;
SharedReg209_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg209_out;
SharedReg210_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg210_out;
Delay60No_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_48_cast <= Delay60No_out;
SharedReg233_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg233_out;
Delay62No4_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_50_cast <= Delay62No4_out;
SharedReg87_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg87_out;
SharedReg173_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg173_out;
SharedReg109_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg109_out;
SharedReg133_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg133_out;
SharedReg144_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg144_out;
SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg58_out;
SharedReg249_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg249_out;
SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg58_out;
SharedReg223_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg223_out;
SharedReg115_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg115_out;
SharedReg184_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg184_out;
SharedReg135_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg135_out;
SharedReg202_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg202_out;
SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg58_out;
   MUX_Product_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg225_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg131_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg101_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg134_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg221_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg63_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg208_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg180_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg230_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg167_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg78_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg59_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg169_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg82_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg84_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg154_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg128_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg76_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg195_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg200_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg212_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg244_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg102_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg113_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg147_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg73_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg188_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg121_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg234_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg92_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg84_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg136_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg67_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg161_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg217_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg88_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => Delay66No2_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg99_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg209_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg210_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => Delay60No_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg233_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => Delay62No4_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg87_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg173_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg109_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg133_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg144_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg249_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg223_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg115_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg74_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg184_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg135_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg202_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg58_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg246_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg240_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg197_out_to_MUX_Product_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product_1_impl_1_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_1_impl_1_out,
                 Y => Delay1No3_out);

Delay1No4_out_to_Product_2_impl_parent_implementedSystem_port_0_cast <= Delay1No4_out;
Delay1No5_out_to_Product_2_impl_parent_implementedSystem_port_1_cast <= Delay1No5_out;
   Product_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product_2_impl_out,
                 X => Delay1No4_out_to_Product_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No5_out_to_Product_2_impl_parent_implementedSystem_port_1_cast);

SharedReg280_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg280_out;
SharedReg312_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg312_out;
SharedReg281_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg281_out;
SharedReg313_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg313_out;
SharedReg282_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg282_out;
SharedReg314_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg314_out;
SharedReg283_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg283_out;
SharedReg315_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg315_out;
SharedReg284_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg284_out;
SharedReg316_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg316_out;
SharedReg288_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg288_out;
SharedReg292_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg292_out;
SharedReg286_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg286_out;
SharedReg261_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg261_out;
SharedReg291_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg291_out;
SharedReg254_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg254_out;
SharedReg285_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg285_out;
SharedReg295_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg295_out;
SharedReg296_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg296_out;
SharedReg263_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg263_out;
SharedReg287_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg287_out;
SharedReg256_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg256_out;
SharedReg299_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg299_out;
SharedReg255_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg255_out;
SharedReg264_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg264_out;
SharedReg267_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg267_out;
SharedReg294_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg294_out;
SharedReg268_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg268_out;
SharedReg300_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg300_out;
SharedReg290_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg290_out;
SharedReg298_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg298_out;
SharedReg258_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg258_out;
SharedReg253_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg253_out;
SharedReg262_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg262_out;
SharedReg265_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg265_out;
SharedReg259_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg259_out;
SharedReg260_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg260_out;
SharedReg297_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg297_out;
SharedReg266_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg266_out;
SharedReg301_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg301_out;
SharedReg302_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg302_out;
SharedReg270_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg270_out;
SharedReg303_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg303_out;
SharedReg271_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg271_out;
SharedReg304_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg304_out;
SharedReg273_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg273_out;
SharedReg305_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg305_out;
SharedReg274_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg274_out;
SharedReg306_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg306_out;
SharedReg289_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg289_out;
SharedReg307_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg307_out;
SharedReg308_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg308_out;
SharedReg269_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg269_out;
SharedReg275_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg275_out;
SharedReg272_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg272_out;
SharedReg276_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg276_out;
SharedReg277_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg277_out;
SharedReg309_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg309_out;
SharedReg310_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg310_out;
SharedReg278_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg278_out;
SharedReg257_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg257_out;
SharedReg293_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg293_out;
SharedReg279_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg279_out;
SharedReg311_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg311_out;
   MUX_Product_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg280_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg312_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg288_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg292_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg286_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg261_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg291_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg254_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg285_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg295_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg296_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg263_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg281_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg287_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg256_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg299_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg255_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg264_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg267_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg294_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg268_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg300_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg290_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg313_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg298_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg258_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg253_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg262_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg265_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg259_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg260_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg297_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg266_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg301_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg282_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg302_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg270_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg303_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg271_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg304_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg273_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg305_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg274_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg306_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg289_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg314_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg307_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg308_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg269_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg275_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg272_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg276_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg277_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg309_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg310_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg278_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg283_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg257_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg293_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg279_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg311_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg315_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg284_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg316_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product_2_impl_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_2_impl_0_out,
                 Y => Delay1No4_out);

SharedReg166_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg166_out;
SharedReg98_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg98_out;
Delay72No_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_3_cast <= Delay72No_out;
SharedReg81_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg81_out;
SharedReg232_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg232_out;
SharedReg216_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg216_out;
SharedReg243_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg243_out;
Delay63No2_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_8_cast <= Delay63No2_out;
SharedReg165_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg165_out;
SharedReg97_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg97_out;
SharedReg65_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg65_out;
SharedReg61_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg61_out;
SharedReg71_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg71_out;
SharedReg101_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg101_out;
SharedReg222_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg222_out;
SharedReg101_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg101_out;
SharedReg107_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg107_out;
SharedReg149_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg149_out;
SharedReg69_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg69_out;
SharedReg178_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg178_out;
SharedReg145_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg145_out;
SharedReg132_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg132_out;
SharedReg113_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg113_out;
SharedReg132_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg132_out;
SharedReg60_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg60_out;
SharedReg103_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg103_out;
SharedReg68_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg68_out;
SharedReg132_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg132_out;
SharedReg75_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg75_out;
SharedReg203_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg203_out;
SharedReg186_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg186_out;
SharedReg219_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg219_out;
SharedReg177_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg177_out;
SharedReg132_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg132_out;
SharedReg104_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg104_out;
SharedReg237_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg237_out;
SharedReg138_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg138_out;
SharedReg152_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg152_out;
SharedReg199_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg199_out;
SharedReg118_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg118_out;
SharedReg90_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg90_out;
SharedReg116_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg116_out;
SharedReg91_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg91_out;
SharedReg119_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg119_out;
SharedReg85_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg85_out;
SharedReg190_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg190_out;
SharedReg170_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg170_out;
SharedReg77_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg77_out;
SharedReg90_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg90_out;
SharedReg65_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg65_out;
SharedReg163_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg163_out;
SharedReg193_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg193_out;
SharedReg187_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg187_out;
SharedReg115_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg115_out;
SharedReg147_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg147_out;
SharedReg206_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg206_out;
SharedReg122_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg122_out;
SharedReg129_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg129_out;
SharedReg93_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg93_out;
SharedReg157_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg157_out;
SharedReg59_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg59_out;
SharedReg63_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_62_cast <= SharedReg63_out;
SharedReg162_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg162_out;
SharedReg172_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg172_out;
   MUX_Product_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg166_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg98_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg65_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg61_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg71_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg101_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg222_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg101_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg107_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg149_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg69_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg178_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => Delay72No_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg145_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg132_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg113_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg132_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg60_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg103_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg68_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg132_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg75_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg203_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg81_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg186_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg219_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg177_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg132_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg104_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg237_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg138_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg152_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg199_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg118_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg232_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg90_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg116_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg91_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg119_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg85_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg190_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg170_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg77_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg90_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg65_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg216_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg163_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg193_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg187_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg115_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg147_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg206_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg122_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg129_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg93_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg157_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg243_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg59_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg63_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg162_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg172_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => Delay63No2_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg165_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg97_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product_2_impl_1_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_2_impl_1_out,
                 Y => Delay1No5_out);

Delay1No6_out_to_Sum1_0_impl_parent_implementedSystem_port_0_cast <= Delay1No6_out;
Delay1No7_out_to_Sum1_0_impl_parent_implementedSystem_port_1_cast <= Delay1No7_out;
   Sum1_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum1_0_impl_out,
                 X => Delay1No6_out_to_Sum1_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No7_out_to_Sum1_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg12_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg12_out;
SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1_out;
SharedReg20_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg20_out;
SharedReg6_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg6_out;
SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1_out;
SharedReg39_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg39_out;
SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1_out;
SharedReg39_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg39_out;
SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg2_out;
SharedReg21_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg21_out;
SharedReg13_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg13_out;
SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg2_out;
SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg2_out;
SharedReg15_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg15_out;
SharedReg34_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg34_out;
SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg2_out;
SharedReg40_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg40_out;
SharedReg14_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg14_out;
SharedReg33_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg33_out;
SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg2_out;
SharedReg40_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg40_out;
SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg2_out;
SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1_out;
SharedReg20_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg20_out;
SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg2_out;
SharedReg21_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg21_out;
SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1_out;
SharedReg17_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg17_out;
SharedReg70_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg70_out;
SharedReg94_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg94_out;
Delay57No2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_33_cast <= Delay57No2_out;
SharedReg140_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg140_out;
SharedReg109_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg109_out;
SharedReg108_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg108_out;
SharedReg224_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg224_out;
SharedReg145_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg145_out;
SharedReg88_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg88_out;
SharedReg165_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg165_out;
SharedReg182_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg182_out;
SharedReg201_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg201_out;
SharedReg72_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg72_out;
SharedReg146_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg146_out;
SharedReg152_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg152_out;
SharedReg209_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg209_out;
SharedReg76_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg76_out;
SharedReg96_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg96_out;
SharedReg130_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg130_out;
SharedReg81_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg81_out;
SharedReg207_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg207_out;
SharedReg228_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg228_out;
SharedReg229_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg229_out;
SharedReg77_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg77_out;
SharedReg83_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg83_out;
SharedReg159_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg159_out;
SharedReg191_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg191_out;
SharedReg84_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg84_out;
SharedReg160_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg160_out;
SharedReg64_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_60_cast <= SharedReg64_out;
SharedReg139_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_61_cast <= SharedReg139_out;
   MUX_Sum1_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_61_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg21_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg13_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg15_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg34_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg40_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg14_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg33_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg40_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg20_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg21_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg17_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg20_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg70_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg94_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => Delay57No2_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg140_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg109_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg108_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg224_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg145_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg88_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg165_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg6_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg182_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg201_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg72_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg146_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg152_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg209_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg76_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg96_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg130_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg81_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg207_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg228_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg229_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg77_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg83_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg159_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg191_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg84_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg160_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg64_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg39_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg139_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_61_cast,
                 iS_7 => SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg39_out_to_MUX_Sum1_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Sum1_0_impl_0_LUT_out,
                 oMux => MUX_Sum1_0_impl_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum1_0_impl_0_out,
                 Y => Delay1No6_out);

SharedReg2_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg11_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg11_out;
SharedReg30_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg30_out;
SharedReg4_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg4_out;
SharedReg4_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg4_out;
SharedReg42_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg42_out;
SharedReg5_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg5_out;
SharedReg43_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg43_out;
SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1_out;
SharedReg20_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg7_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg7_out;
SharedReg14_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg14_out;
SharedReg5_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg5_out;
SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg8_out;
SharedReg27_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg27_out;
SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1_out;
SharedReg39_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg39_out;
SharedReg3_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg3_out;
SharedReg22_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg22_out;
SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1_out;
SharedReg39_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg39_out;
SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1_out;
Delay64No_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_25_cast <= Delay64No_out;
Delay64No1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_26_cast <= Delay64No1_out;
SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1_out;
SharedReg20_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg20_out;
SharedReg2_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg2_out;
SharedReg8_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg8_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg58_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg58_out;
SharedReg61_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg61_out;
SharedReg103_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg103_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg58_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg58_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg58_out;
SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg131_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg58_out;
SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg131_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg58_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg58_out;
SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg131_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg58_out;
SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg131_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg58_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg58_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg58_out;
SharedReg100_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg100_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg58_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg58_out;
SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg131_out;
SharedReg62_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg62_out;
SharedReg62_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg62_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg58_out;
SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg58_out;
SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg131_out;
SharedReg137_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg137_out;
SharedReg179_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg179_out;
SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_60_cast <= SharedReg131_out;
SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_61_cast <= SharedReg131_out;
   MUX_Sum1_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_61_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg2_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg7_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg14_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg5_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg8_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg27_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg39_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg3_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg11_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg22_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg39_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => Delay64No_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => Delay64No1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg20_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg2_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg8_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg30_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg61_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg103_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg4_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg100_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg4_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg62_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg62_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg58_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg137_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg179_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg42_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg131_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_61_cast,
                 iS_7 => SharedReg5_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg43_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1_out_to_MUX_Sum1_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Sum1_0_impl_1_LUT_out,
                 oMux => MUX_Sum1_0_impl_1_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum1_0_impl_1_out,
                 Y => Delay1No7_out);

Delay1No8_out_to_Sum1_1_impl_parent_implementedSystem_port_0_cast <= Delay1No8_out;
Delay1No9_out_to_Sum1_1_impl_parent_implementedSystem_port_1_cast <= Delay1No9_out;
   Sum1_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum1_1_impl_out,
                 X => Delay1No8_out_to_Sum1_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No9_out_to_Sum1_1_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
SharedReg35_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg35_out;
SharedReg50_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg50_out;
SharedReg39_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg39_out;
SharedReg47_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg47_out;
SharedReg40_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg40_out;
SharedReg51_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg51_out;
SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg21_out;
SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg21_out;
SharedReg9_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg9_out;
SharedReg53_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg53_out;
SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg21_out;
SharedReg52_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg52_out;
SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg21_out;
SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg21_out;
SharedReg19_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg19_out;
SharedReg49_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg49_out;
SharedReg18_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg20_out;
SharedReg39_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg39_out;
SharedReg30_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg30_out;
SharedReg55_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg55_out;
SharedReg208_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg208_out;
SharedReg66_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg66_out;
SharedReg86_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg86_out;
SharedReg86_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg86_out;
SharedReg126_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg126_out;
SharedReg76_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg76_out;
SharedReg153_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg153_out;
SharedReg247_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg247_out;
SharedReg155_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg155_out;
SharedReg156_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg156_out;
SharedReg120_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg120_out;
SharedReg160_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg160_out;
   MUX_Sum1_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_34_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg35_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg53_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg52_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg19_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg49_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg18_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg20_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg39_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg50_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg30_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg55_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg208_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg66_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg86_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg86_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg126_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg76_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg153_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg247_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg39_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg155_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg156_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg120_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg160_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_4 => SharedReg47_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg40_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg51_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg21_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg9_out_to_MUX_Sum1_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Sum1_1_impl_0_LUT_out,
                 oMux => MUX_Sum1_1_impl_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum1_1_impl_0_out,
                 Y => Delay1No8_out);

SharedReg25_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg25_out;
SharedReg43_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg43_out;
SharedReg49_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg49_out;
SharedReg39_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg39_out;
SharedReg39_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg39_out;
SharedReg45_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg45_out;
SharedReg20_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg20_out;
SharedReg24_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg24_out;
SharedReg6_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg6_out;
SharedReg46_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg46_out;
SharedReg20_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg46_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg46_out;
SharedReg41_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg41_out;
SharedReg20_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg20_out;
SharedReg2_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg2_out;
SharedReg20_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg20_out;
SharedReg4_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg4_out;
SharedReg27_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg27_out;
SharedReg21_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg21_out;
SharedReg40_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg40_out;
SharedReg46_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg46_out;
SharedReg131_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg131_out;
SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg100_out;
SharedReg131_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg131_out;
SharedReg132_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg132_out;
SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg100_out;
SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg100_out;
SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg100_out;
SharedReg58_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg58_out;
SharedReg131_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg131_out;
SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg100_out;
SharedReg175_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg175_out;
SharedReg197_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg197_out;
SharedReg245_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg245_out;
   MUX_Sum1_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_34_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg43_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg46_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg41_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg20_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg2_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg20_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg4_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg27_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg21_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg40_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg49_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg46_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg131_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg131_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg132_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg58_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg131_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg39_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg100_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg175_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg197_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg245_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_4 => SharedReg39_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg45_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg20_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg24_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg6_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg46_out_to_MUX_Sum1_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Sum1_1_impl_1_LUT_out,
                 oMux => MUX_Sum1_1_impl_1_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum1_1_impl_1_out,
                 Y => Delay1No9_out);

Delay1No10_out_to_Sum1_2_impl_parent_implementedSystem_port_0_cast <= Delay1No10_out;
Delay1No11_out_to_Sum1_2_impl_parent_implementedSystem_port_1_cast <= Delay1No11_out;
   Sum1_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum1_2_impl_out,
                 X => Delay1No10_out_to_Sum1_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No11_out_to_Sum1_2_impl_parent_implementedSystem_port_1_cast);

SharedReg16_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg31_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg31_out;
SharedReg44_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg44_out;
SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg20_out;
SharedReg39_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg39_out;
SharedReg9_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg9_out;
SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg32_out;
SharedReg2_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg2_out;
SharedReg40_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg40_out;
SharedReg21_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg21_out;
SharedReg40_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg40_out;
SharedReg2_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg2_out;
SharedReg40_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg40_out;
SharedReg40_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg40_out;
SharedReg39_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg39_out;
SharedReg11_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg11_out;
SharedReg1_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1_out;
SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg20_out;
SharedReg1_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1_out;
SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg20_out;
SharedReg11_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg11_out;
SharedReg36_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg36_out;
SharedReg67_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg67_out;
SharedReg110_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg110_out;
SharedReg111_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg111_out;
SharedReg171_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg171_out;
SharedReg79_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg79_out;
SharedReg66_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg66_out;
SharedReg183_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg183_out;
SharedReg181_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg181_out;
SharedReg185_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg185_out;
SharedReg168_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg168_out;
SharedReg239_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg239_out;
SharedReg152_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg152_out;
SharedReg149_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg149_out;
SharedReg81_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg81_out;
SharedReg242_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg242_out;
SharedReg250_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg250_out;
SharedReg114_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg114_out;
SharedReg114_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg114_out;
SharedReg150_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg150_out;
SharedReg150_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg150_out;
SharedReg95_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg95_out;
SharedReg215_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg215_out;
SharedReg159_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg159_out;
SharedReg82_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg82_out;
SharedReg82_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg82_out;
SharedReg192_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg192_out;
   MUX_Sum1_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_51_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg16_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg2_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg40_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg21_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg40_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg2_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg40_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg40_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg39_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg11_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg31_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg11_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg36_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg67_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg110_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg111_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg171_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg79_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg44_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg66_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg183_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg181_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg185_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg168_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg239_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg152_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg149_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg81_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg242_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg250_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg114_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg114_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg150_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg150_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg95_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg215_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg159_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg82_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg82_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg192_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_6 => SharedReg39_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg9_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg20_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg32_out_to_MUX_Sum1_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Sum1_2_impl_0_LUT_out,
                 oMux => MUX_Sum1_2_impl_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum1_2_impl_0_out,
                 Y => Delay1No10_out);

SharedReg6_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg6_out;
SharedReg21_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg21_out;
SharedReg24_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg24_out;
SharedReg42_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg42_out;
SharedReg23_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg23_out;
SharedReg1_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1_out;
SharedReg24_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg24_out;
SharedReg26_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg26_out;
SharedReg1_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1_out;
SharedReg33_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg33_out;
SharedReg52_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg52_out;
SharedReg43_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg43_out;
SharedReg20_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg20_out;
SharedReg39_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg39_out;
SharedReg8_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg8_out;
SharedReg39_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg39_out;
Delay64No2_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_17_cast <= Delay64No2_out;
SharedReg2_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg2_out;
SharedReg1_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1_out;
SharedReg39_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg39_out;
SharedReg21_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg21_out;
SharedReg2_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg2_out;
SharedReg21_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg21_out;
SharedReg8_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg8_out;
SharedReg27_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg27_out;
SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg100_out;
SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg131_out;
SharedReg134_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg134_out;
SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg58_out;
SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg58_out;
SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg58_out;
SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg58_out;
SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg131_out;
SharedReg197_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg197_out;
SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg58_out;
SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg131_out;
SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg100_out;
SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg131_out;
SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg58_out;
SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg100_out;
SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg58_out;
SharedReg175_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg175_out;
SharedReg197_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg197_out;
SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg131_out;
SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg131_out;
SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg100_out;
SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg131_out;
SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg100_out;
SharedReg137_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg137_out;
SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg58_out;
SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg100_out;
   MUX_Sum1_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_51_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg6_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg21_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg52_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg43_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg20_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg39_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg8_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg39_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => Delay64No2_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg2_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg39_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg24_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg21_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg2_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg21_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg8_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg27_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg134_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg42_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg197_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg23_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg175_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg197_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg131_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg137_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg58_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg100_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_6 => SharedReg24_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg26_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg33_out_to_MUX_Sum1_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Sum1_2_impl_1_LUT_out,
                 oMux => MUX_Sum1_2_impl_1_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum1_2_impl_1_out,
                 Y => Delay1No11_out);

Delay1No12_out_to_Sum12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No12_out;
Delay1No13_out_to_Sum12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No13_out;
   Sum12_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum12_2_impl_out,
                 X => Delay1No12_out_to_Sum12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No13_out_to_Sum12_2_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
SharedReg54_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg54_out;
SharedReg39_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg39_out;
SharedReg28_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg28_out;
SharedReg28_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg28_out;
SharedReg38_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg38_out;
SharedReg21_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg21_out;
SharedReg10_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg10_out;
SharedReg56_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg56_out;
SharedReg39_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg39_out;
SharedReg49_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg49_out;
SharedReg142_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg142_out;
SharedReg144_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg144_out;
SharedReg79_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg79_out;
SharedReg200_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg200_out;
SharedReg89_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg89_out;
SharedReg214_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg214_out;
SharedReg227_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg227_out;
SharedReg95_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg95_out;
SharedReg155_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg155_out;
   MUX_Sum12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_20_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg54_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg49_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg142_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg144_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg79_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg200_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg89_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg214_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg227_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg95_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg155_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg39_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg28_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg28_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg38_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg21_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg10_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg56_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg39_out_to_MUX_Sum12_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Sum12_2_impl_0_LUT_out,
                 oMux => MUX_Sum12_2_impl_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum12_2_impl_0_out,
                 Y => Delay1No12_out);

SharedReg44_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg44_out;
SharedReg40_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg20_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg25_out;
SharedReg21_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg21_out;
SharedReg20_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg20_out;
SharedReg8_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg8_out;
SharedReg42_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg42_out;
SharedReg40_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg40_out;
SharedReg46_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg46_out;
SharedReg175_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg175_out;
SharedReg58_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg58_out;
SharedReg131_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg131_out;
SharedReg236_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg236_out;
SharedReg100_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg100_out;
SharedReg101_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg101_out;
SharedReg175_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg175_out;
SharedReg58_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg58_out;
SharedReg131_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg131_out;
SharedReg100_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg100_out;
   MUX_Sum12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_20_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg44_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg175_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg58_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg131_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg236_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg100_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg101_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg175_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg58_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg131_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg100_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg20_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg25_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg21_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg20_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg8_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg42_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg40_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg46_out_to_MUX_Sum12_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Sum12_2_impl_1_LUT_out,
                 oMux => MUX_Sum12_2_impl_1_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum12_2_impl_1_out,
                 Y => Delay1No13_out);

Delay1No14_out_to_Sum15_2_impl_parent_implementedSystem_port_0_cast <= Delay1No14_out;
Delay1No15_out_to_Sum15_2_impl_parent_implementedSystem_port_1_cast <= Delay1No15_out;
   Sum15_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum15_2_impl_out,
                 X => Delay1No14_out_to_Sum15_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No15_out_to_Sum15_2_impl_parent_implementedSystem_port_1_cast);

SharedReg40_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg40_out;
SharedReg47_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg47_out;
SharedReg57_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg57_out;
SharedReg48_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg48_out;
SharedReg40_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg40_out;
SharedReg37_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg37_out;
SharedReg89_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg89_out;
SharedReg112_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg112_out;
SharedReg168_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg168_out;
SharedReg130_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg130_out;
SharedReg155_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg155_out;
SharedReg251_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg251_out;
SharedReg64_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg64_out;
   MUX_Sum15_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg40_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg47_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg155_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg251_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg64_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg57_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg48_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg40_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg37_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg89_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg112_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg168_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg130_out_to_MUX_Sum15_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Sum15_2_impl_0_LUT_out,
                 oMux => MUX_Sum15_2_impl_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum15_2_impl_0_out,
                 Y => Delay1No14_out);

SharedReg39_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg39_out;
SharedReg44_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg44_out;
SharedReg40_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg40_out;
SharedReg46_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg46_out;
SharedReg39_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg39_out;
SharedReg23_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg23_out;
SharedReg100_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg100_out;
SharedReg131_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg131_out;
SharedReg175_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg175_out;
SharedReg100_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg100_out;
SharedReg175_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg175_out;
SharedReg105_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg105_out;
SharedReg175_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg175_out;
   MUX_Sum15_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg39_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg44_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg175_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg105_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg175_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg40_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg46_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg39_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg23_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg100_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg131_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg175_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg100_out_to_MUX_Sum15_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Sum15_2_impl_1_LUT_out,
                 oMux => MUX_Sum15_2_impl_1_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum15_2_impl_1_out,
                 Y => Delay1No15_out);

Delay1No16_out_to_Sum2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No16_out;
Delay1No17_out_to_Sum2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No17_out;
   Sum2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum2_2_impl_out,
                 X => Delay1No16_out_to_Sum2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No17_out_to_Sum2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
SharedReg29_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg29_out;
SharedReg39_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg39_out;
SharedReg158_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg158_out;
SharedReg190_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg190_out;
SharedReg80_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg80_out;
   MUX_Sum2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg39_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg158_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg190_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg80_out_to_MUX_Sum2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => MUX_Sum2_2_impl_0_LUT_out,
                 oMux => MUX_Sum2_2_impl_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum2_2_impl_0_out,
                 Y => Delay1No16_out);

SharedReg27_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg27_out;
SharedReg40_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg176_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg176_out;
SharedReg100_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg100_out;
SharedReg218_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg218_out;
SharedReg197_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg197_out;
   MUX_Sum2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg27_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg176_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg100_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg218_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg197_out_to_MUX_Sum2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => MUX_Sum2_2_impl_1_LUT_out,
                 oMux => MUX_Sum2_2_impl_1_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum2_2_impl_1_out,
                 Y => Delay1No17_out);

Delay1No18_out_to_Sum26_1_impl_parent_implementedSystem_port_0_cast <= Delay1No18_out;
Delay1No19_out_to_Sum26_1_impl_parent_implementedSystem_port_1_cast <= Delay1No19_out;
   Sum26_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum26_1_impl_out,
                 X => Delay1No18_out_to_Sum26_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No19_out_to_Sum26_1_impl_parent_implementedSystem_port_1_cast);

SharedReg25_out_to_MUX_Sum26_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg25_out;
SharedReg194_out_to_MUX_Sum26_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg194_out;
SharedReg80_out_to_MUX_Sum26_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg80_out;
   MUX_Sum26_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Sum26_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg194_out_to_MUX_Sum26_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg80_out_to_MUX_Sum26_1_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Sum26_1_impl_0_LUT_out,
                 oMux => MUX_Sum26_1_impl_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum26_1_impl_0_out,
                 Y => Delay1No18_out);

SharedReg23_out_to_MUX_Sum26_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg23_out;
SharedReg100_out_to_MUX_Sum26_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg100_out;
SharedReg197_out_to_MUX_Sum26_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg197_out;
   MUX_Sum26_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg23_out_to_MUX_Sum26_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg100_out_to_MUX_Sum26_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg197_out_to_MUX_Sum26_1_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Sum26_1_impl_1_LUT_out,
                 oMux => MUX_Sum26_1_impl_1_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum26_1_impl_1_out,
                 Y => Delay1No19_out);

Delay1No20_out_to_Sum41_2_impl_parent_implementedSystem_port_0_cast <= Delay1No20_out;
Delay1No21_out_to_Sum41_2_impl_parent_implementedSystem_port_1_cast <= Delay1No21_out;
   Sum41_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum41_2_impl_out,
                 X => Delay1No20_out_to_Sum41_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No21_out_to_Sum41_2_impl_parent_implementedSystem_port_1_cast);

SharedReg30_out_to_MUX_Sum41_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg30_out;
SharedReg155_out_to_MUX_Sum41_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg155_out;
   MUX_Sum41_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg30_out_to_MUX_Sum41_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg155_out_to_MUX_Sum41_2_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Sum41_2_impl_0_LUT_out,
                 oMux => MUX_Sum41_2_impl_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum41_2_impl_0_out,
                 Y => Delay1No20_out);

SharedReg27_out_to_MUX_Sum41_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg27_out;
SharedReg197_out_to_MUX_Sum41_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg197_out;
   MUX_Sum41_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg27_out_to_MUX_Sum41_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg197_out_to_MUX_Sum41_2_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Sum41_2_impl_1_LUT_out,
                 oMux => MUX_Sum41_2_impl_1_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum41_2_impl_1_out,
                 Y => Delay1No21_out);

Delay1No22_out_to_Sum42_2_impl_parent_implementedSystem_port_0_cast <= Delay1No22_out;
Delay1No23_out_to_Sum42_2_impl_parent_implementedSystem_port_1_cast <= Delay1No23_out;
   Sum42_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum42_2_impl_out,
                 X => Delay1No22_out_to_Sum42_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No23_out_to_Sum42_2_impl_parent_implementedSystem_port_1_cast);

SharedReg72_out_to_MUX_Sum42_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg117_out_to_MUX_Sum42_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Sum42_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_Sum42_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Sum42_2_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Sum42_2_impl_0_LUT_out,
                 oMux => MUX_Sum42_2_impl_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum42_2_impl_0_out,
                 Y => Delay1No22_out);

SharedReg175_out_to_MUX_Sum42_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg175_out;
SharedReg218_out_to_MUX_Sum42_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg218_out;
   MUX_Sum42_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg175_out_to_MUX_Sum42_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg218_out_to_MUX_Sum42_2_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Sum42_2_impl_1_LUT_out,
                 oMux => MUX_Sum42_2_impl_1_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum42_2_impl_1_out,
                 Y => Delay1No23_out);
   a_0_impl_instance: Constant_float_8_23_0_617123672897668340553423149685841053724_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a_0_impl_out);
   a1_0_impl_instance: Constant_float_8_23_0_631862801488796588245122620719484984875_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a1_0_impl_out);
   a10_0_impl_instance: Constant_float_8_23_1_436934552725145586293820088030770421028_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a10_0_impl_out);
   a11_0_impl_instance: Constant_float_8_23_1_561088850170149200380365073215216398239_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a11_0_impl_out);
   a12_0_impl_instance: Constant_float_8_23_1_67381401040949318037576176720904186368_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a12_0_impl_out);
   a13_0_impl_instance: Constant_float_8_23_1_767419732788928943278961014584638178349_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a13_0_impl_out);
   a14_0_impl_instance: Constant_float_8_23_1_83466961525726479642628419242100790143_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a14_0_impl_out);
   a15_0_impl_instance: Constant_float_8_23_1_869869533302351394254969818575773388147_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a15_0_impl_out);
   a2_0_impl_instance: Constant_float_8_23_0_663686724095854829741369940165895968676_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a2_0_impl_out);
   a3_0_impl_instance: Constant_float_8_23_0_712333225863809871292176012502750381827_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a3_0_impl_out);
   a4_0_impl_instance: Constant_float_8_23_0_777424256340159325340266605053329840302_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a4_0_impl_out);
   a5_0_impl_instance: Constant_float_8_23_0_858338451424324633265428019512910395861_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a5_0_impl_out);
   a6_0_impl_instance: Constant_float_8_23_0_95403875322976861017565397560247220099_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a6_0_impl_out);
   a7_0_impl_instance: Constant_float_8_23_1_062858000783881262663044253713451325893_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a7_0_impl_out);
   a8_0_impl_instance: Constant_float_8_23_1_182256984960216694702239692560397088528_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a8_0_impl_out);
   a9_0_impl_instance: Constant_float_8_23_1_308589307952890523623068474989850074053_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => a9_0_impl_out);
   b_0_impl_instance: Constant_float_8_23_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => b_0_impl_out);
   c_0_impl_instance: Constant_float_8_23_n0_99584180311675085661704542872030287981_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c_0_impl_out);
   c1_0_impl_instance: Constant_float_8_23_n0_987534845729581944873132215434452518821_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c1_0_impl_out);
   c10_0_impl_instance: Constant_float_8_23_n0_906979034015293006376623452524654567242_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c10_0_impl_out);
   c11_0_impl_instance: Constant_float_8_23_n0_898568629504465254953515795932617038488_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c11_0_impl_out);
   c12_0_impl_instance: Constant_float_8_23_n0_891139475905879052675118145998567342758_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c12_0_impl_out);
   c13_0_impl_instance: Constant_float_8_23_n0_885091234632599865861379839770961552858_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c13_0_impl_out);
   c14_0_impl_instance: Constant_float_8_23_n0_880803415623673480183697392931208014488_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c14_0_impl_out);
   c15_0_impl_instance: Constant_float_8_23_n0_878576235602384070233483726042322814465_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c15_0_impl_out);
   c2_0_impl_instance: Constant_float_8_23_n0_979173278459382512295405831537209451199_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c2_0_impl_out);
   c3_0_impl_instance: Constant_float_8_23_n0_970685163049390786760284299816703423858_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c3_0_impl_out);
   c4_0_impl_instance: Constant_float_8_23_n0_962013487567665803723571116279345005751_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c4_0_impl_out);
   c5_0_impl_instance: Constant_float_8_23_n0_95312319664069156122110371143207885325_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c5_0_impl_out);
   c6_0_impl_instance: Constant_float_8_23_n0_944010225685960935315677033941028639674_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c6_0_impl_out);
   c7_0_impl_instance: Constant_float_8_23_n0_934712586109242460352675152535084635019_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c7_0_impl_out);
   c8_0_impl_instance: Constant_float_8_23_n0_925322845902050161726037913467735052109_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c8_0_impl_out);
   c9_0_impl_instance: Constant_float_8_23_n0_916000226493365876656582713621901348233_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => c9_0_impl_out);
   d_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => d_0_impl_out);
   Out2_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Out2_0_IEEE,
                 X => Delay1No24_out);
Out2_0 <= Out2_0_IEEE;

SharedReg58_out_to_MUX_Out2_0_0_parent_implementedSystem_port_1_cast <= SharedReg58_out;
SharedReg175_out_to_MUX_Out2_0_0_parent_implementedSystem_port_2_cast <= SharedReg175_out;
SharedReg100_out_to_MUX_Out2_0_0_parent_implementedSystem_port_3_cast <= SharedReg100_out;
   MUX_Out2_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg58_out_to_MUX_Out2_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg175_out_to_MUX_Out2_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg100_out_to_MUX_Out2_0_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Out2_0_0_LUT_out,
                 oMux => MUX_Out2_0_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Out2_0_0_out,
                 Y => Delay1No24_out);

   Delay64No_instance: Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=37 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg19_out,
                 Y => Delay64No_out);

   Delay64No1_instance: Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=37 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => Delay64No1_out);

   Delay64No2_instance: Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=37 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => Delay64No2_out);

   Delay57No2_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => Delay57No2_out);

   Delay60No_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => Delay60No_out);

   Delay63No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => Delay63No2_out);

   Delay63No3_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => Delay63No3_out);

   Delay62No4_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => Delay62No4_out);

   Delay72No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => Delay72No_out);

   Delay71No1_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => Delay71No1_out);

   Delay67No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => Delay67No1_out);

   Delay66No2_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => Delay66No2_out);

   MUX_Sum1_0_impl_0_LUT_instance: GenericLut_LUTData_MUX_Sum1_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum1_0_impl_0_LUT_out);

   MUX_Sum1_0_impl_1_LUT_instance: GenericLut_LUTData_MUX_Sum1_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum1_0_impl_1_LUT_out);

   MUX_Sum1_1_impl_0_LUT_instance: GenericLut_LUTData_MUX_Sum1_1_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum1_1_impl_0_LUT_out);

   MUX_Sum1_1_impl_1_LUT_instance: GenericLut_LUTData_MUX_Sum1_1_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum1_1_impl_1_LUT_out);

   MUX_Sum1_2_impl_0_LUT_instance: GenericLut_LUTData_MUX_Sum1_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum1_2_impl_0_LUT_out);

   MUX_Sum1_2_impl_1_LUT_instance: GenericLut_LUTData_MUX_Sum1_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum1_2_impl_1_LUT_out);

   MUX_Sum12_2_impl_0_LUT_instance: GenericLut_LUTData_MUX_Sum12_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum12_2_impl_0_LUT_out);

   MUX_Sum12_2_impl_1_LUT_instance: GenericLut_LUTData_MUX_Sum12_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum12_2_impl_1_LUT_out);

   MUX_Sum15_2_impl_0_LUT_instance: GenericLut_LUTData_MUX_Sum15_2_impl_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum15_2_impl_0_LUT_out);

   MUX_Sum15_2_impl_1_LUT_instance: GenericLut_LUTData_MUX_Sum15_2_impl_1_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum15_2_impl_1_LUT_out);

   MUX_Sum2_2_impl_0_LUT_instance: GenericLut_LUTData_MUX_Sum2_2_impl_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum2_2_impl_0_LUT_out);

   MUX_Sum2_2_impl_1_LUT_instance: GenericLut_LUTData_MUX_Sum2_2_impl_1_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum2_2_impl_1_LUT_out);

   MUX_Sum26_1_impl_0_LUT_instance: GenericLut_LUTData_MUX_Sum26_1_impl_0_LUT_wIn_6_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum26_1_impl_0_LUT_out);

   MUX_Sum26_1_impl_1_LUT_instance: GenericLut_LUTData_MUX_Sum26_1_impl_1_LUT_wIn_6_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum26_1_impl_1_LUT_out);

   MUX_Sum41_2_impl_0_LUT_instance: GenericLut_LUTData_MUX_Sum41_2_impl_0_LUT_wIn_6_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum41_2_impl_0_LUT_out);

   MUX_Sum41_2_impl_1_LUT_instance: GenericLut_LUTData_MUX_Sum41_2_impl_1_LUT_wIn_6_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum41_2_impl_1_LUT_out);

   MUX_Sum42_2_impl_0_LUT_instance: GenericLut_LUTData_MUX_Sum42_2_impl_0_LUT_wIn_6_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum42_2_impl_0_LUT_out);

   MUX_Sum42_2_impl_1_LUT_instance: GenericLut_LUTData_MUX_Sum42_2_impl_1_LUT_wIn_6_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Sum42_2_impl_1_LUT_out);

   MUX_Out2_0_0_LUT_instance: GenericLut_LUTData_MUX_Out2_0_0_LUT_wIn_6_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Out2_0_0_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=68 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => In2_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product_0_impl_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg2_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg3_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg4_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg6_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg7_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg8_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg9_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg10_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg11_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg12_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg13_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg14_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg15_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg16_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg17_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg18_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product_1_impl_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg20_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg21_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg22_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg23_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg24_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg25_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg26_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg27_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg28_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg29_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg30_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg31_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product_2_impl_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum1_0_impl_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum1_1_impl_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum1_2_impl_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum12_2_impl_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum15_2_impl_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum2_2_impl_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum26_1_impl_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum41_2_impl_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum42_2_impl_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a_0_impl_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_100_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=100 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a1_0_impl_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_684_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=684 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a10_0_impl_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_746_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=746 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a11_0_impl_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_849_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=849 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a12_0_impl_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_948_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=948 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a13_0_impl_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_1016_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1016 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a14_0_impl_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_1081_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1081 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a15_0_impl_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_162_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=162 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a2_0_impl_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_246_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=246 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a3_0_impl_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_296_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=296 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a4_0_impl_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_365_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=365 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a5_0_impl_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_439_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=439 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a6_0_impl_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_507_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=507 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a7_0_impl_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_558_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=558 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a8_0_impl_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_624_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=624 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => a9_0_impl_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_73_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=73 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => b_0_impl_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_75_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=75 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=55 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_70_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=70 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=65 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=67 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=67 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_130_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=130 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=37 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c_0_impl_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=97 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c1_0_impl_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_681_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=681 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c10_0_impl_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_735_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=735 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c11_0_impl_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_838_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=838 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c12_0_impl_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_946_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=946 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c13_0_impl_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_995_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=995 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c14_0_impl_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_1056_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1056 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c15_0_impl_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_146_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=146 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c2_0_impl_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_239_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=239 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c3_0_impl_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_294_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=294 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c4_0_impl_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_359_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=359 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c5_0_impl_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_442_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=442 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c6_0_impl_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_499_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=499 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c7_0_impl_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_555_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=555 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c8_0_impl_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_625_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=625 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => c9_0_impl_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=60 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => d_0_impl_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=65 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=65 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_70_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=70 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=65 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=69 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_130_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=130 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => SharedReg316_out);
end architecture;

