--------------------------------------------------------------------------------
--                         ModuloCounter_7_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_7_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of ModuloCounter_7_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(2 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 6 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_2_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(0 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0",
         iS_1 when "1",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid2164070_RightShifter
--                (RightShifter_24_by_max_26_F250_uid2164072)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2164070_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2164070_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid2164075
--                  (IntAdderAlternative_27_f250_uid2164079)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid2164075 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid2164075 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid2164082
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid2164082 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid2164082 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid2164085
--                   (IntAdderClassical_34_f250_uid2164087)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid2164085 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid2164085 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid2164070
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2164070 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2164070 is
   component FPAdd_8_23_uid2164070_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid2164075 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid2164082 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid2164085 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid2164070_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid2164075  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid2164082  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid2164085  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid2164070 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid2164070  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_7_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_7_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_7_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
         iS_5 when "101",
         iS_6 when "110",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2165127
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2165127 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2165127 is
signal XX_m2165128 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m2165128 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m2165128 <= X ;
   YY_m2165128 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid2165131
--                   (IntAdderClassical_33_f500_uid2165133)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid2165131 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid2165131 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2165127 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid2165131 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2165127  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid2165131  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid2165258_RightShifter
--                (RightShifter_24_by_max_26_F250_uid2165260)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2165258_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2165258_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid2165263
--                  (IntAdderAlternative_27_f250_uid2165267)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid2165263 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid2165263 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid2165270
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid2165270 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid2165270 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid2165273
--                   (IntAdderClassical_34_f250_uid2165275)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid2165273 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid2165273 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid2165258
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2165258 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2165258 is
   component FPAdd_8_23_uid2165258_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid2165263 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid2165270 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid2165273 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid2165258_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid2165263  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid2165270  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid2165273  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid2165258 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid2165258  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_6_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_6_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_6_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
         iS_5 when "101",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_0_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "1" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "1" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "1" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "1" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "1" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "1" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "1" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "1" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "1" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "1" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "1" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "1" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "1" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "1" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "1" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "1" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "1" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "1" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "1" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "1" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "1" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "1" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "1" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "1" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "1" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "1" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "1" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "1" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "1" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "1" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "1" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "0" when "011",
      "1" when "100",
      "0" when "101",
      "0" when "110",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product331_1_impl_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product331_1_impl_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product331_1_impl_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "101" when "000",
      "001" when "001",
      "010" when "010",
      "000" when "011",
      "000" when "100",
      "011" when "101",
      "100" when "110",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product331_1_impl_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product331_1_impl_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product331_1_impl_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Product331_1_impl_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_Product331_1_impl_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product331_1_impl_1_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product331_1_impl_1_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product331_1_impl_1_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "010" when "000",
      "011" when "001",
      "100" when "010",
      "000" when "011",
      "101" when "100",
      "000" when "101",
      "001" when "110",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product331_1_impl_1_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product331_1_impl_1_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product331_1_impl_1_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Product331_1_impl_1_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_Product331_1_impl_1_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      Y <= s15;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      Y <= s17;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          x0_re_0 : in std_logic_vector(31 downto 0);
          x0_im_0 : in std_logic_vector(31 downto 0);
          x1_re_0 : in std_logic_vector(31 downto 0);
          x1_im_0 : in std_logic_vector(31 downto 0);
          x2_re_0 : in std_logic_vector(31 downto 0);
          x2_im_0 : in std_logic_vector(31 downto 0);
          x3_re_0 : in std_logic_vector(31 downto 0);
          x3_im_0 : in std_logic_vector(31 downto 0);
          x4_re_0 : in std_logic_vector(31 downto 0);
          x4_im_0 : in std_logic_vector(31 downto 0);
          x5_re_0 : in std_logic_vector(31 downto 0);
          x5_im_0 : in std_logic_vector(31 downto 0);
          x6_re_0 : in std_logic_vector(31 downto 0);
          x6_im_0 : in std_logic_vector(31 downto 0);
          x7_re_0 : in std_logic_vector(31 downto 0);
          x7_im_0 : in std_logic_vector(31 downto 0);
          x8_re_0 : in std_logic_vector(31 downto 0);
          x8_im_0 : in std_logic_vector(31 downto 0);
          x9_re_0 : in std_logic_vector(31 downto 0);
          x9_im_0 : in std_logic_vector(31 downto 0);
          x10_re_0 : in std_logic_vector(31 downto 0);
          x10_im_0 : in std_logic_vector(31 downto 0);
          x11_re_0 : in std_logic_vector(31 downto 0);
          x11_im_0 : in std_logic_vector(31 downto 0);
          x12_re_0 : in std_logic_vector(31 downto 0);
          x12_im_0 : in std_logic_vector(31 downto 0);
          x13_re_0 : in std_logic_vector(31 downto 0);
          x13_im_0 : in std_logic_vector(31 downto 0);
          x14_re_0 : in std_logic_vector(31 downto 0);
          x14_im_0 : in std_logic_vector(31 downto 0);
          x15_re_0 : in std_logic_vector(31 downto 0);
          x15_im_0 : in std_logic_vector(31 downto 0);
          y0_re_0 : out std_logic_vector(31 downto 0);
          y0_im_0 : out std_logic_vector(31 downto 0);
          y1_re_0 : out std_logic_vector(31 downto 0);
          y1_im_0 : out std_logic_vector(31 downto 0);
          y2_re_0 : out std_logic_vector(31 downto 0);
          y2_im_0 : out std_logic_vector(31 downto 0);
          y3_re_0 : out std_logic_vector(31 downto 0);
          y3_im_0 : out std_logic_vector(31 downto 0);
          y4_re_0 : out std_logic_vector(31 downto 0);
          y4_im_0 : out std_logic_vector(31 downto 0);
          y5_re_0 : out std_logic_vector(31 downto 0);
          y5_im_0 : out std_logic_vector(31 downto 0);
          y6_re_0 : out std_logic_vector(31 downto 0);
          y6_im_0 : out std_logic_vector(31 downto 0);
          y7_re_0 : out std_logic_vector(31 downto 0);
          y7_im_0 : out std_logic_vector(31 downto 0);
          y8_re_0 : out std_logic_vector(31 downto 0);
          y8_im_0 : out std_logic_vector(31 downto 0);
          y9_re_0 : out std_logic_vector(31 downto 0);
          y9_im_0 : out std_logic_vector(31 downto 0);
          y10_re_0 : out std_logic_vector(31 downto 0);
          y10_im_0 : out std_logic_vector(31 downto 0);
          y11_re_0 : out std_logic_vector(31 downto 0);
          y11_im_0 : out std_logic_vector(31 downto 0);
          y12_re_0 : out std_logic_vector(31 downto 0);
          y12_im_0 : out std_logic_vector(31 downto 0);
          y13_re_0 : out std_logic_vector(31 downto 0);
          y13_im_0 : out std_logic_vector(31 downto 0);
          y14_re_0 : out std_logic_vector(31 downto 0);
          y14_im_0 : out std_logic_vector(31 downto 0);
          y15_re_0 : out std_logic_vector(31 downto 0);
          y15_im_0 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_7_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(2 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_2_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(0 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_7_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_6_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product331_1_impl_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product331_1_impl_1_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount71_out : std_logic_vector(2 downto 0) := (others => '0');
signal x0_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add16_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add117_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add117_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add117_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add117_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add117_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add117_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add120_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add120_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add120_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add120_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add120_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add120_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add36_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add36_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add36_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add36_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add36_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add36_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add127_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add127_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add127_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add127_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add127_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add127_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add38_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add38_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add38_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add38_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add38_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add38_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add128_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add128_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add129_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add129_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add40_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add40_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add130_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add130_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product13_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product25_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product25_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product25_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product25_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product25_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product25_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product35_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product35_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product35_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product35_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product35_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product35_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract6_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product9_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product16_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product16_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product16_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product16_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product16_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product36_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product36_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product36_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product36_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product36_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product36_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract7_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract23_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract23_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product124_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product124_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product323_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product323_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product324_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product324_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product324_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product324_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product324_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product324_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product325_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product325_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product325_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product226_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product226_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product130_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product130_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product130_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product329_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product329_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product329_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product329_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product329_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product329_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract30_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract30_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product132_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product132_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product132_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product132_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product132_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product132_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product331_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product331_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product331_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product331_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product331_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product331_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract42_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract42_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract44_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract44_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract45_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract45_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract45_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract45_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract45_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract45_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract46_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract46_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract57_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract57_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract57_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract57_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract57_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract57_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract117_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract117_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract117_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract117_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract117_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract117_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract61_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract61_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract61_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract61_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract61_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract61_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract121_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract121_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract121_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract121_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract121_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract121_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant14_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant15_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant8_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant17_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y0_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y1_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y1_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y2_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y2_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y3_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y3_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y4_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y4_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y5_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y5_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y6_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y6_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y7_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y7_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y8_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y8_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y9_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y9_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y10_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y10_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y11_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y11_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y12_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y12_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y13_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y13_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y14_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y14_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y15_re_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_y15_im_0_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product331_1_impl_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Product331_1_impl_1_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No1_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No10_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No11_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Add16_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Add16_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Add16_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Add16_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Add9_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Add9_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Add9_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Add9_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Add18_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Add18_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No8_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Add18_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Add18_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No19_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No9_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Add117_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Add117_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No4_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Add117_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Add117_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No5_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Add120_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Add120_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Add120_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Add120_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Add36_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Add36_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No32_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No34_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Add36_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Add36_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No33_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No35_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Add127_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Add127_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No84_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No8_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Add127_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Add127_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No9_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No41_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Add38_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Add38_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No56_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No46_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Add38_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Add38_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No57_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Add128_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Add128_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No26_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No44_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No68_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Add128_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Add128_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No27_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No47_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Add129_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Add129_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No36_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Add129_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Add129_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No37_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Add40_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Add40_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Add40_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Add40_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Add130_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Add130_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Add130_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Add130_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Product11_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Product11_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Product11_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Product11_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Product5_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Product5_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Product5_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Product5_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Subtract3_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Subtract3_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No30_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No12_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No6_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Subtract3_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Subtract3_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No31_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No7_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No13_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Product13_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Product13_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Product13_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Product13_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Product25_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Product25_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Product25_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Product25_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Product35_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Product35_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out_to_Product35_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out_to_Product35_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out_to_Subtract6_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out_to_Subtract6_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No66_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No86_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No28_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No10_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out_to_Subtract6_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out_to_Subtract6_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No67_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No29_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No11_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No87_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out_to_Product9_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out_to_Product9_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out_to_Product9_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out_to_Product9_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out_to_Product16_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out_to_Product16_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out_to_Product16_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out_to_Product16_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out_to_Product26_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out_to_Product26_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out_to_Product26_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out_to_Product26_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out_to_Product36_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out_to_Product36_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out_to_Product36_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out_to_Product36_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out_to_Subtract7_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out_to_Subtract7_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out_to_Subtract7_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out_to_Subtract7_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out_to_Product18_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out_to_Product18_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out_to_Product18_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out_to_Product18_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out_to_Product28_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out_to_Product28_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out_to_Product28_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out_to_Product28_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out_to_Subtract9_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out_to_Subtract9_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No42_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No48_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out_to_Subtract9_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out_to_Subtract9_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No43_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No49_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out_to_Product221_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out_to_Product221_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out_to_Product221_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out_to_Product221_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out_to_Product321_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out_to_Product321_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out_to_Product321_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out_to_Product321_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out_to_Subtract23_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out_to_Subtract23_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No22_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out_to_Subtract23_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out_to_Subtract23_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No23_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out_to_Product124_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out_to_Product124_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out_to_Product124_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out_to_Product124_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out_to_Product323_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out_to_Product323_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out_to_Product323_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out_to_Product323_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out_to_Product324_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out_to_Product324_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out_to_Product324_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out_to_Product324_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out_to_Product325_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out_to_Product325_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out_to_Product55_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out_to_Product55_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out_to_Product226_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out_to_Product226_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out_to_Product226_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out_to_Product226_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out_to_Product130_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out_to_Product130_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out_to_Product329_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out_to_Product329_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out_to_Product329_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out_to_Product329_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out_to_Subtract30_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out_to_Subtract30_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No32_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out_to_Subtract30_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out_to_Subtract30_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No33_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out_to_Product132_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out_to_Product132_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out_to_Product132_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out_to_Product132_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out_to_Product331_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out_to_Product331_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No8_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out_to_Product331_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out_to_Product331_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No9_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out_to_Subtract42_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out_to_Subtract42_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out_to_Subtract42_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out_to_Subtract42_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out_to_Subtract44_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out_to_Subtract44_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out_to_Subtract44_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out_to_Subtract44_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out_to_Subtract45_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out_to_Subtract45_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out_to_Subtract45_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out_to_Subtract45_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out_to_Subtract46_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out_to_Subtract46_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out_to_Subtract46_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out_to_Subtract46_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out_to_Subtract57_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out_to_Subtract57_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out_to_Subtract57_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out_to_Subtract57_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out_to_Subtract117_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out_to_Subtract117_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out_to_Subtract117_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out_to_Subtract117_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out_to_Subtract61_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out_to_Subtract61_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out_to_Subtract61_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out_to_Subtract61_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out_to_Subtract121_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out_to_Subtract121_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out_to_Subtract121_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out_to_Subtract121_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount71_instance: ModuloCounter_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount71_out);
x0_re_0_IEEE <= x0_re_0;
   x0_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_re_0_out,
                 X => x0_re_0_IEEE);
x0_im_0_IEEE <= x0_im_0;
   x0_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_im_0_out,
                 X => x0_im_0_IEEE);
x1_re_0_IEEE <= x1_re_0;
   x1_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_re_0_out,
                 X => x1_re_0_IEEE);
x1_im_0_IEEE <= x1_im_0;
   x1_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_im_0_out,
                 X => x1_im_0_IEEE);
x2_re_0_IEEE <= x2_re_0;
   x2_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_re_0_out,
                 X => x2_re_0_IEEE);
x2_im_0_IEEE <= x2_im_0;
   x2_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_im_0_out,
                 X => x2_im_0_IEEE);
x3_re_0_IEEE <= x3_re_0;
   x3_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_re_0_out,
                 X => x3_re_0_IEEE);
x3_im_0_IEEE <= x3_im_0;
   x3_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_im_0_out,
                 X => x3_im_0_IEEE);
x4_re_0_IEEE <= x4_re_0;
   x4_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_re_0_out,
                 X => x4_re_0_IEEE);
x4_im_0_IEEE <= x4_im_0;
   x4_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_im_0_out,
                 X => x4_im_0_IEEE);
x5_re_0_IEEE <= x5_re_0;
   x5_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_re_0_out,
                 X => x5_re_0_IEEE);
x5_im_0_IEEE <= x5_im_0;
   x5_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_im_0_out,
                 X => x5_im_0_IEEE);
x6_re_0_IEEE <= x6_re_0;
   x6_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_re_0_out,
                 X => x6_re_0_IEEE);
x6_im_0_IEEE <= x6_im_0;
   x6_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_im_0_out,
                 X => x6_im_0_IEEE);
x7_re_0_IEEE <= x7_re_0;
   x7_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_re_0_out,
                 X => x7_re_0_IEEE);
x7_im_0_IEEE <= x7_im_0;
   x7_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_im_0_out,
                 X => x7_im_0_IEEE);
x8_re_0_IEEE <= x8_re_0;
   x8_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_re_0_out,
                 X => x8_re_0_IEEE);
x8_im_0_IEEE <= x8_im_0;
   x8_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_im_0_out,
                 X => x8_im_0_IEEE);
x9_re_0_IEEE <= x9_re_0;
   x9_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_re_0_out,
                 X => x9_re_0_IEEE);
x9_im_0_IEEE <= x9_im_0;
   x9_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_im_0_out,
                 X => x9_im_0_IEEE);
x10_re_0_IEEE <= x10_re_0;
   x10_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_re_0_out,
                 X => x10_re_0_IEEE);
x10_im_0_IEEE <= x10_im_0;
   x10_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_im_0_out,
                 X => x10_im_0_IEEE);
x11_re_0_IEEE <= x11_re_0;
   x11_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_re_0_out,
                 X => x11_re_0_IEEE);
x11_im_0_IEEE <= x11_im_0;
   x11_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_im_0_out,
                 X => x11_im_0_IEEE);
x12_re_0_IEEE <= x12_re_0;
   x12_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_re_0_out,
                 X => x12_re_0_IEEE);
x12_im_0_IEEE <= x12_im_0;
   x12_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_im_0_out,
                 X => x12_im_0_IEEE);
x13_re_0_IEEE <= x13_re_0;
   x13_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_re_0_out,
                 X => x13_re_0_IEEE);
x13_im_0_IEEE <= x13_im_0;
   x13_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_im_0_out,
                 X => x13_im_0_IEEE);
x14_re_0_IEEE <= x14_re_0;
   x14_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_re_0_out,
                 X => x14_re_0_IEEE);
x14_im_0_IEEE <= x14_im_0;
   x14_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_im_0_out,
                 X => x14_im_0_IEEE);
x15_re_0_IEEE <= x15_re_0;
   x15_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_re_0_out,
                 X => x15_re_0_IEEE);
x15_im_0_IEEE <= x15_im_0;
   x15_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_im_0_out,
                 X => x15_im_0_IEEE);
   y0_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_re_0_IEEE,
                 X => Delay1No_out);
y0_re_0 <= y0_re_0_IEEE;

SharedReg38_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg38_out;
SharedReg41_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg41_out;
   MUX_y0_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg38_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg41_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y0_re_0_0_LUT_out,
                 oMux => MUX_y0_re_0_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_re_0_0_out,
                 Y => Delay1No_out);
   y0_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_im_0_IEEE,
                 X => Delay1No1_out);
y0_im_0 <= y0_im_0_IEEE;

SharedReg44_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg44_out;
SharedReg49_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg49_out;
   MUX_y0_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg44_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg49_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y0_im_0_0_LUT_out,
                 oMux => MUX_y0_im_0_0_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_im_0_0_out,
                 Y => Delay1No1_out);
   y1_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_re_0_IEEE,
                 X => Delay1No2_out);
y1_re_0 <= y1_re_0_IEEE;

SharedReg60_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg63_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg63_out;
   MUX_y1_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg63_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y1_re_0_0_LUT_out,
                 oMux => MUX_y1_re_0_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_re_0_0_out,
                 Y => Delay1No2_out);
   y1_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_im_0_IEEE,
                 X => Delay1No3_out);
y1_im_0 <= y1_im_0_IEEE;

SharedReg66_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg66_out;
SharedReg69_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg69_out;
   MUX_y1_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg66_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg69_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y1_im_0_0_LUT_out,
                 oMux => MUX_y1_im_0_0_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_im_0_0_out,
                 Y => Delay1No3_out);
   y2_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_re_0_IEEE,
                 X => Delay1No4_out);
y2_re_0 <= y2_re_0_IEEE;

SharedReg78_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg78_out;
SharedReg81_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg81_out;
   MUX_y2_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg78_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg81_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y2_re_0_0_LUT_out,
                 oMux => MUX_y2_re_0_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_re_0_0_out,
                 Y => Delay1No4_out);
   y2_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_im_0_IEEE,
                 X => Delay1No5_out);
y2_im_0 <= y2_im_0_IEEE;

SharedReg84_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg84_out;
SharedReg87_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg87_out;
   MUX_y2_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg84_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg87_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y2_im_0_0_LUT_out,
                 oMux => MUX_y2_im_0_0_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_im_0_0_out,
                 Y => Delay1No5_out);
   y3_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_re_0_IEEE,
                 X => Delay1No6_out);
y3_re_0 <= y3_re_0_IEEE;

SharedReg38_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg38_out;
SharedReg41_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg41_out;
   MUX_y3_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg38_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg41_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y3_re_0_0_LUT_out,
                 oMux => MUX_y3_re_0_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_re_0_0_out,
                 Y => Delay1No6_out);
   y3_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_im_0_IEEE,
                 X => Delay1No7_out);
y3_im_0 <= y3_im_0_IEEE;

SharedReg44_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg44_out;
SharedReg49_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg49_out;
   MUX_y3_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg44_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg49_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y3_im_0_0_LUT_out,
                 oMux => MUX_y3_im_0_0_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_im_0_0_out,
                 Y => Delay1No7_out);
   y4_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_re_0_IEEE,
                 X => Delay1No8_out);
y4_re_0 <= y4_re_0_IEEE;

SharedReg57_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg57_out;
SharedReg54_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg54_out;
   MUX_y4_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg57_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg54_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y4_re_0_0_LUT_out,
                 oMux => MUX_y4_re_0_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_re_0_0_out,
                 Y => Delay1No8_out);
   y4_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_im_0_IEEE,
                 X => Delay1No9_out);
y4_im_0 <= y4_im_0_IEEE;

SharedReg60_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg63_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg63_out;
   MUX_y4_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg63_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y4_im_0_0_LUT_out,
                 oMux => MUX_y4_im_0_0_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_im_0_0_out,
                 Y => Delay1No9_out);
   y5_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_re_0_IEEE,
                 X => Delay1No10_out);
y5_re_0 <= y5_re_0_IEEE;

SharedReg78_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg78_out;
SharedReg81_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg81_out;
   MUX_y5_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg78_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg81_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y5_re_0_0_LUT_out,
                 oMux => MUX_y5_re_0_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_re_0_0_out,
                 Y => Delay1No10_out);
   y5_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_im_0_IEEE,
                 X => Delay1No11_out);
y5_im_0 <= y5_im_0_IEEE;

SharedReg84_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg84_out;
SharedReg87_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg87_out;
   MUX_y5_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg84_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg87_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y5_im_0_0_LUT_out,
                 oMux => MUX_y5_im_0_0_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_im_0_0_out,
                 Y => Delay1No11_out);
   y6_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_re_0_IEEE,
                 X => Delay1No12_out);
y6_re_0 <= y6_re_0_IEEE;

SharedReg66_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg66_out;
SharedReg69_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg69_out;
   MUX_y6_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg66_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg69_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y6_re_0_0_LUT_out,
                 oMux => MUX_y6_re_0_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_re_0_0_out,
                 Y => Delay1No12_out);
   y6_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_im_0_IEEE,
                 X => Delay1No13_out);
y6_im_0 <= y6_im_0_IEEE;

SharedReg72_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg75_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg75_out;
   MUX_y6_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg75_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y6_im_0_0_LUT_out,
                 oMux => MUX_y6_im_0_0_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_im_0_0_out,
                 Y => Delay1No13_out);
   y7_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_re_0_IEEE,
                 X => Delay1No14_out);
y7_re_0 <= y7_re_0_IEEE;

SharedReg90_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg90_out;
SharedReg93_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg93_out;
   MUX_y7_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg90_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg93_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y7_re_0_0_LUT_out,
                 oMux => MUX_y7_re_0_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_re_0_0_out,
                 Y => Delay1No14_out);
   y7_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_im_0_IEEE,
                 X => Delay1No15_out);
y7_im_0 <= y7_im_0_IEEE;

SharedReg54_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg54_out;
SharedReg57_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg57_out;
   MUX_y7_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg54_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg57_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y7_im_0_0_LUT_out,
                 oMux => MUX_y7_im_0_0_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_im_0_0_out,
                 Y => Delay1No15_out);
   y8_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_re_0_IEEE,
                 X => Delay1No16_out);
y8_re_0 <= y8_re_0_IEEE;

SharedReg380_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg380_out;
SharedReg383_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg383_out;
   MUX_y8_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg380_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg383_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y8_re_0_0_LUT_out,
                 oMux => MUX_y8_re_0_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_re_0_0_out,
                 Y => Delay1No16_out);
   y8_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_im_0_IEEE,
                 X => Delay1No17_out);
y8_im_0 <= y8_im_0_IEEE;

SharedReg386_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg386_out;
SharedReg388_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg388_out;
   MUX_y8_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg386_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg388_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y8_im_0_0_LUT_out,
                 oMux => MUX_y8_im_0_0_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_im_0_0_out,
                 Y => Delay1No17_out);
   y9_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_re_0_IEEE,
                 X => Delay1No18_out);
y9_re_0 <= y9_re_0_IEEE;

SharedReg372_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg372_out;
SharedReg376_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg376_out;
   MUX_y9_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg372_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg376_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y9_re_0_0_LUT_out,
                 oMux => MUX_y9_re_0_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_re_0_0_out,
                 Y => Delay1No18_out);
   y9_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_im_0_IEEE,
                 X => Delay1No19_out);
y9_im_0 <= y9_im_0_IEEE;

SharedReg380_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg380_out;
SharedReg383_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg383_out;
   MUX_y9_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg380_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg383_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y9_im_0_0_LUT_out,
                 oMux => MUX_y9_im_0_0_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_im_0_0_out,
                 Y => Delay1No19_out);
   y10_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_re_0_IEEE,
                 X => Delay1No20_out);
y10_re_0 <= y10_re_0_IEEE;

SharedReg358_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg358_out;
SharedReg362_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg362_out;
   MUX_y10_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg358_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg362_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y10_re_0_0_LUT_out,
                 oMux => MUX_y10_re_0_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_re_0_0_out,
                 Y => Delay1No20_out);
   y10_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_im_0_IEEE,
                 X => Delay1No21_out);
y10_im_0 <= y10_im_0_IEEE;

SharedReg290_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg290_out;
SharedReg296_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg296_out;
   MUX_y10_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg290_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg296_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y10_im_0_0_LUT_out,
                 oMux => MUX_y10_im_0_0_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_im_0_0_out,
                 Y => Delay1No21_out);
   y11_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_re_0_IEEE,
                 X => Delay1No22_out);
y11_re_0 <= y11_re_0_IEEE;

SharedReg350_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg350_out;
SharedReg354_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg354_out;
   MUX_y11_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg350_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg354_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y11_re_0_0_LUT_out,
                 oMux => MUX_y11_re_0_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_re_0_0_out,
                 Y => Delay1No22_out);
   y11_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_im_0_IEEE,
                 X => Delay1No23_out);
y11_im_0 <= y11_im_0_IEEE;

SharedReg366_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg366_out;
SharedReg369_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg369_out;
   MUX_y11_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg366_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg369_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y11_im_0_0_LUT_out,
                 oMux => MUX_y11_im_0_0_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_im_0_0_out,
                 Y => Delay1No23_out);
   y12_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_re_0_IEEE,
                 X => Delay1No24_out);
y12_re_0 <= y12_re_0_IEEE;

SharedReg390_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg391_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg391_out;
   MUX_y12_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y12_re_0_0_LUT_out,
                 oMux => MUX_y12_re_0_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_re_0_0_out,
                 Y => Delay1No24_out);
   y12_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_im_0_IEEE,
                 X => Delay1No25_out);
y12_im_0 <= y12_im_0_IEEE;

SharedReg326_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg326_out;
SharedReg331_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg331_out;
   MUX_y12_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg326_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg331_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y12_im_0_0_LUT_out,
                 oMux => MUX_y12_im_0_0_out);

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_im_0_0_out,
                 Y => Delay1No25_out);
   y13_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_re_0_IEEE,
                 X => Delay1No26_out);
y13_re_0 <= y13_re_0_IEEE;

SharedReg386_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg386_out;
SharedReg388_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg388_out;
   MUX_y13_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg386_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg388_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y13_re_0_0_LUT_out,
                 oMux => MUX_y13_re_0_0_out);

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_re_0_0_out,
                 Y => Delay1No26_out);
   y13_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_im_0_IEEE,
                 X => Delay1No27_out);
y13_im_0 <= y13_im_0_IEEE;

SharedReg390_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg391_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg391_out;
   MUX_y13_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y13_im_0_0_LUT_out,
                 oMux => MUX_y13_im_0_0_out);

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_im_0_0_out,
                 Y => Delay1No27_out);
   y14_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_re_0_IEEE,
                 X => Delay1No28_out);
y14_re_0 <= y14_re_0_IEEE;

SharedReg358_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg358_out;
SharedReg362_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg362_out;
   MUX_y14_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg358_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg362_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y14_re_0_0_LUT_out,
                 oMux => MUX_y14_re_0_0_out);

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_re_0_0_out,
                 Y => Delay1No28_out);
   y14_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_im_0_IEEE,
                 X => Delay1No29_out);
y14_im_0 <= y14_im_0_IEEE;

SharedReg326_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg326_out;
SharedReg331_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg331_out;
   MUX_y14_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg326_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg331_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y14_im_0_0_LUT_out,
                 oMux => MUX_y14_im_0_0_out);

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_im_0_0_out,
                 Y => Delay1No29_out);
   y15_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_re_0_IEEE,
                 X => Delay1No30_out);
y15_re_0 <= y15_re_0_IEEE;

SharedReg386_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg386_out;
SharedReg388_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg388_out;
   MUX_y15_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg386_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg388_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y15_re_0_0_LUT_out,
                 oMux => MUX_y15_re_0_0_out);

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_re_0_0_out,
                 Y => Delay1No30_out);
   y15_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_im_0_IEEE,
                 X => Delay1No31_out);
y15_im_0 <= y15_im_0_IEEE;

SharedReg390_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg391_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg391_out;
   MUX_y15_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_y15_im_0_0_LUT_out,
                 oMux => MUX_y15_im_0_0_out);

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_im_0_0_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Add2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_0_impl_out,
                 X => Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg215_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg215_out;
SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg136_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg136_out;
SharedReg254_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg254_out;
SharedReg173_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg173_out;
SharedReg92_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg92_out;
SharedReg174_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg174_out;
   MUX_Add2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg215_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg136_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg254_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg173_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg92_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg174_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add2_0_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_0_out,
                 Y => Delay1No32_out);

SharedReg171_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg171_out;
SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg146_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg146_out;
SharedReg341_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg341_out;
SharedReg366_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg366_out;
SharedReg72_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg72_out;
SharedReg190_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg190_out;
   MUX_Add2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg171_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg146_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg341_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg366_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg72_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg190_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add2_0_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Add2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_1_impl_out,
                 X => Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg258_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg258_out;
SharedReg177_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg177_out;
SharedReg95_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg95_out;
SharedReg178_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg178_out;
SharedReg218_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg218_out;
SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg_out;
SharedReg141_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg141_out;
   MUX_Add2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg258_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg177_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg95_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg178_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg218_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg141_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add2_1_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_0_out,
                 Y => Delay1No34_out);

SharedReg346_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg346_out;
SharedReg369_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg369_out;
SharedReg75_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg75_out;
SharedReg194_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg194_out;
SharedReg175_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg175_out;
SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg16_out;
SharedReg151_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg151_out;
   MUX_Add2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg346_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg369_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg75_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg194_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg151_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add2_1_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Add11_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_0_impl_out,
                 X => Delay1No36_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast);

SharedReg96_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg96_out;
SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg270_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg270_out;
SharedReg255_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg255_out;
SharedReg188_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg188_out;
SharedReg99_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg99_out;
SharedReg189_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg189_out;
   MUX_Add11_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg96_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg270_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg255_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg188_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg99_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg189_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add11_0_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_0_out,
                 Y => Delay1No36_out);

SharedReg104_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg104_out;
SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg233_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg233_out;
SharedReg344_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg344_out;
SharedReg171_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg171_out;
SharedReg146_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg146_out;
SharedReg257_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg257_out;
   MUX_Add11_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg104_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg233_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg344_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg171_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg146_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg257_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add11_0_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Add11_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_1_impl_out,
                 X => Delay1No38_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast);

SharedReg259_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg259_out;
SharedReg192_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg192_out;
SharedReg103_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg103_out;
SharedReg193_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg193_out;
SharedReg100_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg100_out;
SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1_out;
SharedReg274_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg274_out;
   MUX_Add11_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg259_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg192_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg103_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg193_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg100_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg274_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add11_1_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_0_out,
                 Y => Delay1No38_out);

SharedReg349_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg349_out;
SharedReg175_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg175_out;
SharedReg151_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg151_out;
SharedReg261_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg261_out;
SharedReg109_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg109_out;
SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg17_out;
SharedReg236_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg236_out;
   MUX_Add11_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg349_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg175_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg151_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg261_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg109_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg236_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add11_1_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Add3_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_0_impl_out,
                 X => Delay1No40_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast);

SharedReg187_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg187_out;
SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg2_out;
SharedReg137_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg137_out;
SharedReg126_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg126_out;
Delay7No_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast <= Delay7No_out;
SharedReg217_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg217_out;
SharedReg91_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg91_out;
   MUX_Add3_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg187_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg137_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg126_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay7No_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg217_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg91_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add3_0_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_0_impl_0_out,
                 Y => Delay1No40_out);

SharedReg233_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg233_out;
SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg96_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg96_out;
SharedReg139_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg139_out;
SharedReg107_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg107_out;
SharedReg215_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg215_out;
SharedReg108_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg108_out;
   MUX_Add3_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg233_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg96_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg139_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg107_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg215_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg108_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add3_0_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_0_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Add3_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_1_impl_out,
                 X => Delay1No42_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast);

SharedReg132_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg132_out;
Delay7No1_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast <= Delay7No1_out;
SharedReg220_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg220_out;
SharedReg94_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg94_out;
SharedReg191_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg191_out;
SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg2_out;
SharedReg142_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg142_out;
   MUX_Add3_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg132_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay7No1_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg220_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg94_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg191_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg142_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add3_1_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_1_impl_0_out,
                 Y => Delay1No42_out);

SharedReg144_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg144_out;
SharedReg112_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg218_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg218_out;
SharedReg113_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg113_out;
SharedReg236_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg236_out;
SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg18_out;
SharedReg100_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg100_out;
   MUX_Add3_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg144_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg218_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg113_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg236_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg100_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add3_1_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_1_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Add12_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_0_impl_out,
                 X => Delay1No44_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg86_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg86_out;
SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg291_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg291_out;
SharedReg149_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg149_out;
SharedReg235_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg235_out;
SharedReg216_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg216_out;
SharedReg271_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg271_out;
   MUX_Add12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg86_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg291_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg149_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg235_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg216_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg271_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add12_0_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_0_impl_0_out,
                 Y => Delay1No44_out);

SharedReg114_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg114_out;
SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg254_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg254_out;
Delay7No10_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast <= Delay7No10_out;
SharedReg292_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg292_out;
SharedReg187_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg187_out;
SharedReg330_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg330_out;
   MUX_Add12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg114_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg254_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay7No10_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg292_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg187_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg330_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add12_0_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_0_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Add12_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_1_impl_out,
                 X => Delay1No46_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg154_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg154_out;
SharedReg238_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg238_out;
SharedReg219_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg219_out;
SharedReg275_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg275_out;
SharedReg89_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg89_out;
SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg3_out;
SharedReg297_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg297_out;
   MUX_Add12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg154_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg238_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg219_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg275_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg89_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg297_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add12_1_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_1_impl_0_out,
                 Y => Delay1No46_out);

Delay7No11_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast <= Delay7No11_out;
SharedReg298_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg298_out;
SharedReg191_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg191_out;
SharedReg335_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg335_out;
SharedReg119_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg119_out;
SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg19_out;
SharedReg258_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg258_out;
   MUX_Add12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay7No11_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg298_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg191_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg335_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg119_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg258_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add12_1_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_1_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Add16_0_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Add16_0_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Add16_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add16_0_impl_out,
                 X => Delay1No48_out_to_Add16_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Add16_0_impl_parent_implementedSystem_port_1_cast);

SharedReg254_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg254_out;
SharedReg4_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg4_out;
SharedReg147_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg147_out;
SharedReg172_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg172_out;
SharedReg117_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg117_out;
SharedReg91_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg91_out;
SharedReg116_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg116_out;
   MUX_Add16_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg254_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg4_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg147_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg172_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg117_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg91_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg116_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add16_0_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_0_impl_0_out,
                 Y => Delay1No48_out);

SharedReg256_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg256_out;
SharedReg20_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg104_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg104_out;
SharedReg269_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg269_out;
SharedReg126_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg126_out;
SharedReg90_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg90_out;
SharedReg140_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg140_out;
   MUX_Add16_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg256_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg104_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg269_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg126_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg90_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg140_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add16_0_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_0_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Add16_1_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Add16_1_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Add16_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add16_1_impl_out,
                 X => Delay1No50_out_to_Add16_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Add16_1_impl_parent_implementedSystem_port_1_cast);

SharedReg176_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg176_out;
SharedReg122_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg122_out;
SharedReg94_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg94_out;
SharedReg121_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg121_out;
SharedReg258_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg258_out;
SharedReg4_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg4_out;
SharedReg152_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg152_out;
   MUX_Add16_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg176_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg122_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg94_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg121_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg258_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg4_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg152_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add16_1_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_1_impl_0_out,
                 Y => Delay1No50_out);

SharedReg273_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg273_out;
SharedReg132_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg132_out;
SharedReg93_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg93_out;
SharedReg145_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg145_out;
SharedReg260_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg260_out;
SharedReg20_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg20_out;
SharedReg109_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg109_out;
   MUX_Add16_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg273_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg132_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg93_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg145_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg260_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg20_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg109_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add16_1_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_1_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Add9_0_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Add9_0_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Add9_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_0_impl_out,
                 X => Delay1No52_out_to_Add9_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Add9_0_impl_parent_implementedSystem_port_1_cast);

SharedReg124_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg124_out;
SharedReg5_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg215_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg215_out;
SharedReg85_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg85_out;
SharedReg172_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg172_out;
SharedReg234_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg234_out;
SharedReg234_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg234_out;
   MUX_Add9_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg124_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg215_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg85_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg172_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg234_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg234_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add9_0_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_0_impl_0_out,
                 Y => Delay1No52_out);

SharedReg107_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg107_out;
SharedReg21_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg21_out;
SharedReg269_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg269_out;
SharedReg136_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg136_out;
SharedReg215_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg215_out;
SharedReg233_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg233_out;
SharedReg295_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg295_out;
   MUX_Add9_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg107_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg21_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg269_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg136_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg215_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg233_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg295_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add9_0_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_0_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Add9_1_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Add9_1_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Add9_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_1_impl_out,
                 X => Delay1No54_out_to_Add9_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Add9_1_impl_parent_implementedSystem_port_1_cast);

SharedReg88_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg88_out;
SharedReg176_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg176_out;
SharedReg237_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg237_out;
SharedReg237_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg237_out;
SharedReg130_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg130_out;
SharedReg5_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg5_out;
SharedReg218_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg218_out;
   MUX_Add9_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg88_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg176_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg237_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg237_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg130_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg5_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg218_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add9_1_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_1_impl_0_out,
                 Y => Delay1No54_out);

SharedReg141_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg141_out;
SharedReg218_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg218_out;
SharedReg236_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg236_out;
SharedReg301_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg301_out;
SharedReg112_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg112_out;
SharedReg21_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg21_out;
SharedReg273_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg273_out;
   MUX_Add9_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg141_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg218_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg236_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg301_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg112_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg21_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg273_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add9_1_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_1_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Add18_0_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Add18_0_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Add18_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_0_impl_out,
                 X => Delay1No56_out_to_Add18_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Add18_0_impl_parent_implementedSystem_port_1_cast);

SharedReg223_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg223_out;
SharedReg12_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg12_out;
SharedReg90_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg90_out;
SharedReg188_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg188_out;
SharedReg97_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg97_out;
SharedReg116_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg116_out;
SharedReg98_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg98_out;
   MUX_Add18_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg223_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg90_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg188_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg97_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg116_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg98_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add18_0_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_0_impl_0_out,
                 Y => Delay1No56_out);

SharedReg156_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg156_out;
SharedReg28_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg28_out;
SharedReg114_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg114_out;
SharedReg358_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg358_out;
SharedReg78_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg78_out;
SharedReg96_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg96_out;
Delay16No8_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_7_cast <= Delay16No8_out;
   MUX_Add18_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg156_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg28_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg114_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg358_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg78_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg96_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay16No8_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add18_0_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_0_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Add18_1_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Add18_1_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Add18_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_1_impl_out,
                 X => Delay1No58_out_to_Add18_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Add18_1_impl_parent_implementedSystem_port_1_cast);

SharedReg192_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg192_out;
SharedReg101_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg101_out;
SharedReg121_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg121_out;
SharedReg102_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg102_out;
Delay5No19_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_5_cast <= Delay5No19_out;
SharedReg12_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg12_out;
SharedReg93_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg93_out;
   MUX_Add18_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg192_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg101_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg121_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg102_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay5No19_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg12_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg93_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add18_1_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_1_impl_0_out,
                 Y => Delay1No58_out);

SharedReg362_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg362_out;
SharedReg81_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg81_out;
SharedReg100_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg100_out;
Delay16No9_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_4_cast <= Delay16No9_out;
SharedReg169_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg169_out;
SharedReg28_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg28_out;
SharedReg119_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg119_out;
   MUX_Add18_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg362_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg81_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg100_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay16No9_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg169_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg28_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg119_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add18_1_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_1_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Add117_0_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Add117_0_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Add117_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add117_0_impl_out,
                 X => Delay1No60_out_to_Add117_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Add117_0_impl_parent_implementedSystem_port_1_cast);

SharedReg163_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg163_out;
SharedReg6_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg6_out;
SharedReg271_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg271_out;
SharedReg86_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg86_out;
SharedReg105_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg105_out;
SharedReg329_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg329_out;
SharedReg210_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg210_out;
   MUX_Add117_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg163_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg6_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg271_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg86_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg105_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg329_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg210_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add117_0_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add117_0_impl_0_out,
                 Y => Delay1No60_out);

SharedReg179_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg179_out;
SharedReg22_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg22_out;
SharedReg294_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg294_out;
SharedReg146_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg146_out;
SharedReg84_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg84_out;
Delay15No4_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_6_cast <= Delay15No4_out;
SharedReg179_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg179_out;
   MUX_Add117_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg179_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg22_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg294_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg146_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg84_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay15No4_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg179_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add117_0_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add117_0_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Add117_1_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Add117_1_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Add117_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add117_1_impl_out,
                 X => Delay1No62_out_to_Add117_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Add117_1_impl_parent_implementedSystem_port_1_cast);

SharedReg89_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg89_out;
SharedReg110_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg110_out;
SharedReg334_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg334_out;
SharedReg213_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg213_out;
SharedReg166_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg166_out;
SharedReg6_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg6_out;
SharedReg275_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg275_out;
   MUX_Add117_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg89_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg110_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg334_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg213_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg166_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg6_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg275_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add117_1_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add117_1_impl_0_out,
                 Y => Delay1No62_out);

SharedReg151_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg151_out;
SharedReg87_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg87_out;
Delay15No5_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_3_cast <= Delay15No5_out;
SharedReg181_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg181_out;
SharedReg185_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg185_out;
SharedReg22_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg22_out;
SharedReg300_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg300_out;
   MUX_Add117_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg151_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg87_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay15No5_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg181_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg185_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg22_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg300_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add117_1_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add117_1_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Add120_0_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Add120_0_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Add120_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add120_0_impl_out,
                 X => Delay1No64_out_to_Add120_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Add120_0_impl_parent_implementedSystem_port_1_cast);

SharedReg184_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg184_out;
SharedReg7_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg7_out;
SharedReg138_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg138_out;
SharedReg167_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg167_out;
SharedReg163_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg163_out;
SharedReg126_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg126_out;
SharedReg221_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg221_out;
   MUX_Add120_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg184_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg138_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg167_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg163_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg126_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg221_out_to_MUX_Add120_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add120_0_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add120_0_impl_0_out,
                 Y => Delay1No64_out);

SharedReg195_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg195_out;
SharedReg23_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg23_out;
SharedReg128_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg128_out;
SharedReg179_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg179_out;
SharedReg167_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg167_out;
SharedReg118_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg118_out;
SharedReg320_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg320_out;
   MUX_Add120_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg195_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg23_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg128_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg179_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg167_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg118_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg320_out_to_MUX_Add120_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add120_0_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add120_0_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Add120_1_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Add120_1_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Add120_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add120_1_impl_out,
                 X => Delay1No66_out_to_Add120_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Add120_1_impl_parent_implementedSystem_port_1_cast);

SharedReg169_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg169_out;
SharedReg166_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg166_out;
SharedReg132_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg132_out;
SharedReg224_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg224_out;
SharedReg186_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg186_out;
SharedReg7_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg7_out;
SharedReg143_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg143_out;
   MUX_Add120_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg169_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg166_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg132_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg224_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg186_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg7_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg143_out_to_MUX_Add120_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add120_1_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add120_1_impl_0_out,
                 Y => Delay1No66_out);

SharedReg181_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg181_out;
SharedReg169_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg169_out;
SharedReg123_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg123_out;
SharedReg322_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg322_out;
SharedReg202_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg202_out;
SharedReg23_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg23_out;
SharedReg134_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg134_out;
   MUX_Add120_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg181_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg169_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg123_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg322_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg202_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg23_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg134_out_to_MUX_Add120_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add120_1_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add120_1_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Add36_0_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Add36_0_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Add36_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add36_0_impl_out,
                 X => Delay1No68_out_to_Add36_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Add36_0_impl_parent_implementedSystem_port_1_cast);

SharedReg251_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg251_out;
SharedReg8_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
SharedReg292_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg292_out;
SharedReg200_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg200_out;
SharedReg195_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg195_out;
SharedReg156_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg156_out;
Delay5No32_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_7_cast <= Delay5No32_out;
   MUX_Add36_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg251_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg292_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg200_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg195_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg156_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay5No32_out_to_MUX_Add36_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add36_0_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add36_0_impl_0_out,
                 Y => Delay1No68_out);

SharedReg227_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg227_out;
SharedReg24_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg353_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg353_out;
SharedReg204_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg204_out;
SharedReg200_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg200_out;
SharedReg167_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg167_out;
Delay5No34_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_7_cast <= Delay5No34_out;
   MUX_Add36_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg227_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg353_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg204_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg200_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg167_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay5No34_out_to_MUX_Add36_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add36_0_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add36_0_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Add36_1_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Add36_1_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Add36_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add36_1_impl_out,
                 X => Delay1No70_out_to_Add36_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Add36_1_impl_parent_implementedSystem_port_1_cast);

SharedReg202_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg202_out;
SharedReg197_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg197_out;
SharedReg159_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg159_out;
Delay5No33_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_4_cast <= Delay5No33_out;
SharedReg253_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg253_out;
SharedReg8_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg8_out;
SharedReg298_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg298_out;
   MUX_Add36_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg202_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg197_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg159_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay5No33_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg253_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg8_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg298_out_to_MUX_Add36_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add36_1_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add36_1_impl_0_out,
                 Y => Delay1No70_out);

SharedReg207_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg207_out;
SharedReg202_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg202_out;
SharedReg169_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg169_out;
Delay5No35_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_4_cast <= Delay5No35_out;
SharedReg241_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg241_out;
SharedReg24_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg24_out;
SharedReg357_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg357_out;
   MUX_Add36_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg207_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg202_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg169_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay5No35_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg241_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg24_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg357_out_to_MUX_Add36_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add36_1_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add36_1_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Add127_0_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Add127_0_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Add127_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add127_0_impl_out,
                 X => Delay1No72_out_to_Add127_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Add127_0_impl_parent_implementedSystem_port_1_cast);

Delay3No84_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_1_cast <= Delay3No84_out;
SharedReg9_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg9_out;
SharedReg180_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg180_out;
SharedReg250_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg250_out;
SharedReg209_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg209_out;
SharedReg195_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg195_out;
Delay6No8_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_7_cast <= Delay6No8_out;
   MUX_Add127_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No84_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg9_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg180_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg250_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg209_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg195_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay6No8_out_to_MUX_Add127_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add127_0_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add127_0_impl_0_out,
                 Y => Delay1No72_out);

SharedReg244_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg244_out;
SharedReg25_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg25_out;
SharedReg184_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg184_out;
SharedReg262_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg262_out;
SharedReg221_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg221_out;
SharedReg200_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg200_out;
SharedReg229_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg229_out;
   MUX_Add127_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg244_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg25_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg184_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg262_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg221_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg200_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg229_out_to_MUX_Add127_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add127_0_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add127_0_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Add127_1_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Add127_1_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Add127_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add127_1_impl_out,
                 X => Delay1No74_out_to_Add127_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Add127_1_impl_parent_implementedSystem_port_1_cast);

SharedReg252_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg252_out;
SharedReg212_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg212_out;
SharedReg197_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg197_out;
Delay6No9_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_4_cast <= Delay6No9_out;
SharedReg306_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg306_out;
SharedReg9_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg9_out;
SharedReg186_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg186_out;
   MUX_Add127_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg252_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg212_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg197_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay6No9_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg306_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg9_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg186_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add127_1_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add127_1_impl_0_out,
                 Y => Delay1No74_out);

SharedReg264_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg264_out;
SharedReg224_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg224_out;
SharedReg202_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg202_out;
Delay5No41_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_4_cast <= Delay5No41_out;
SharedReg249_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg249_out;
SharedReg25_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg198_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg198_out;
   MUX_Add127_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg264_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg224_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg202_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay5No41_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg249_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg25_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg198_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add127_1_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add127_1_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Add38_0_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Add38_0_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Add38_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add38_0_impl_out,
                 X => Delay1No76_out_to_Add38_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Add38_0_impl_parent_implementedSystem_port_1_cast);

SharedReg204_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg204_out;
SharedReg10_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg10_out;
SharedReg205_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg205_out;
Delay3No56_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_4_cast <= Delay3No56_out;
SharedReg244_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg244_out;
SharedReg239_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg239_out;
SharedReg244_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg244_out;
   MUX_Add38_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg204_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg205_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay3No56_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg244_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg239_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg244_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add38_0_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add38_0_impl_0_out,
                 Y => Delay1No76_out);

SharedReg209_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg209_out;
SharedReg26_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg26_out;
Delay3No46_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_3_cast <= Delay3No46_out;
SharedReg164_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg164_out;
SharedReg248_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg248_out;
SharedReg244_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg244_out;
SharedReg248_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg248_out;
   MUX_Add38_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg209_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg26_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No46_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg164_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg248_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg244_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg248_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add38_0_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add38_0_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Add38_1_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Add38_1_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Add38_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add38_1_impl_out,
                 X => Delay1No78_out_to_Add38_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Add38_1_impl_parent_implementedSystem_port_1_cast);

Delay3No57_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_1_cast <= Delay3No57_out;
SharedReg246_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg246_out;
SharedReg241_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg241_out;
SharedReg246_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg246_out;
SharedReg212_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg212_out;
SharedReg10_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg10_out;
SharedReg213_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg213_out;
   MUX_Add38_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No57_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg246_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg241_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg246_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg212_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg10_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg213_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add38_1_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add38_1_impl_0_out,
                 Y => Delay1No78_out);

SharedReg161_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg161_out;
SharedReg249_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg249_out;
SharedReg246_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg246_out;
SharedReg249_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg249_out;
SharedReg224_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg224_out;
SharedReg26_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg26_out;
SharedReg199_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg199_out;
   MUX_Add38_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg161_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg249_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg246_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg249_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg224_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg26_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg199_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add38_1_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add38_1_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Add128_0_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Add128_0_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Add128_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add128_0_impl_out,
                 X => Delay1No80_out_to_Add128_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Add128_0_impl_parent_implementedSystem_port_1_cast);

SharedReg262_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg262_out;
SharedReg11_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg11_out;
SharedReg303_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg303_out;
Delay5No26_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_4_cast <= Delay5No26_out;
SharedReg240_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg240_out;
SharedReg265_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg265_out;
Delay5No44_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_7_cast <= Delay5No44_out;
   MUX_Add128_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg262_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg11_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg303_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay5No26_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg240_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg265_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay5No44_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add128_0_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_0_impl_0_out,
                 Y => Delay1No80_out);

SharedReg265_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg265_out;
SharedReg27_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg27_out;
SharedReg308_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg308_out;
Delay3No68_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_4_cast <= Delay3No68_out;
SharedReg265_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg265_out;
SharedReg277_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg277_out;
SharedReg280_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg280_out;
   MUX_Add128_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg265_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg308_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay3No68_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg265_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg277_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg280_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add128_0_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_0_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Add128_1_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Add128_1_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Add128_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add128_1_impl_out,
                 X => Delay1No82_out_to_Add128_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Add128_1_impl_parent_implementedSystem_port_1_cast);

Delay5No27_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_1_cast <= Delay5No27_out;
SharedReg242_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg242_out;
SharedReg267_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg267_out;
SharedReg284_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg284_out;
SharedReg267_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg267_out;
SharedReg11_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg11_out;
SharedReg310_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg310_out;
   MUX_Add128_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No27_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg242_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg267_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg284_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg267_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg11_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg310_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add128_1_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_1_impl_0_out,
                 Y => Delay1No82_out);

SharedReg253_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg253_out;
SharedReg267_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg267_out;
SharedReg281_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg281_out;
Delay5No47_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_4_cast <= Delay5No47_out;
SharedReg281_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg281_out;
SharedReg27_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg27_out;
SharedReg314_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg314_out;
   MUX_Add128_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg253_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg267_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg281_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay5No47_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg281_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg27_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg314_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add128_1_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_1_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Add129_0_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Add129_0_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Add129_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add129_0_impl_out,
                 X => Delay1No84_out_to_Add129_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Add129_0_impl_parent_implementedSystem_port_1_cast);

SharedReg302_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg302_out;
SharedReg13_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg244_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg244_out;
SharedReg184_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg184_out;
SharedReg263_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg263_out;
Delay5No36_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_6_cast <= Delay5No36_out;
SharedReg265_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg265_out;
   MUX_Add129_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg302_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg244_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg184_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg263_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay5No36_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg265_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add129_0_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_0_impl_0_out,
                 Y => Delay1No84_out);

SharedReg307_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg307_out;
SharedReg29_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg29_out;
SharedReg248_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg248_out;
SharedReg196_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg196_out;
SharedReg266_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg266_out;
SharedReg211_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg211_out;
SharedReg277_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg277_out;
   MUX_Add129_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg307_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg248_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg196_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg266_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg211_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg277_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add129_0_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_0_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Add129_1_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Add129_1_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Add129_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add129_1_impl_out,
                 X => Delay1No86_out_to_Add129_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Add129_1_impl_parent_implementedSystem_port_1_cast);

SharedReg198_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg198_out;
SharedReg268_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg268_out;
Delay5No37_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_3_cast <= Delay5No37_out;
SharedReg267_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg267_out;
SharedReg309_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg309_out;
SharedReg13_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg13_out;
SharedReg249_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg249_out;
   MUX_Add129_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg198_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg268_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay5No37_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg267_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg309_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg13_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg249_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add129_1_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_1_impl_0_out,
                 Y => Delay1No86_out);

SharedReg203_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg203_out;
SharedReg283_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg283_out;
SharedReg226_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg226_out;
SharedReg281_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg281_out;
SharedReg313_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg313_out;
SharedReg29_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg29_out;
SharedReg252_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg252_out;
   MUX_Add129_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg203_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg283_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg226_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg281_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg313_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg29_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg252_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add129_1_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_1_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Add40_0_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Add40_0_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Add40_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add40_0_impl_out,
                 X => Delay1No88_out_to_Add40_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Add40_0_impl_parent_implementedSystem_port_1_cast);

SharedReg319_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg319_out;
SharedReg14_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg14_out;
SharedReg307_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg307_out;
SharedReg307_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg307_out;
SharedReg285_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg285_out;
SharedReg308_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg308_out;
SharedReg307_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg307_out;
   MUX_Add40_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg319_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg14_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg307_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg307_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg285_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg308_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg307_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add40_0_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_0_impl_0_out,
                 Y => Delay1No88_out);

SharedReg324_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg324_out;
SharedReg30_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg30_out;
SharedReg311_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg311_out;
SharedReg311_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg311_out;
SharedReg302_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg302_out;
SharedReg336_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg336_out;
SharedReg311_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg311_out;
   MUX_Add40_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg324_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg311_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg311_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg302_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg336_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg311_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add40_0_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_0_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Add40_1_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Add40_1_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Add40_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add40_1_impl_out,
                 X => Delay1No90_out_to_Add40_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Add40_1_impl_parent_implementedSystem_port_1_cast);

SharedReg309_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg309_out;
SharedReg288_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg288_out;
SharedReg310_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg310_out;
SharedReg309_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg309_out;
SharedReg323_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg323_out;
SharedReg14_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg14_out;
SharedReg313_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg313_out;
   MUX_Add40_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg309_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg288_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg310_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg309_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg323_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg14_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg313_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add40_1_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_1_impl_0_out,
                 Y => Delay1No90_out);

SharedReg313_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg313_out;
SharedReg304_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg304_out;
SharedReg325_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg325_out;
SharedReg313_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg313_out;
SharedReg325_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg325_out;
SharedReg30_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg30_out;
SharedReg315_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg315_out;
   MUX_Add40_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg313_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg304_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg325_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg313_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg325_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg30_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg315_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add40_1_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_1_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Add130_0_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Add130_0_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Add130_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add130_0_impl_out,
                 X => Delay1No92_out_to_Add130_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Add130_0_impl_parent_implementedSystem_port_1_cast);

SharedReg280_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg280_out;
SharedReg15_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg324_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg324_out;
SharedReg324_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg324_out;
SharedReg336_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg336_out;
SharedReg318_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg318_out;
SharedReg324_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg324_out;
   MUX_Add130_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg280_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg324_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg324_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg336_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg318_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg324_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add130_0_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_0_impl_0_out,
                 Y => Delay1No92_out);

SharedReg338_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg338_out;
SharedReg31_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg31_out;
SharedReg336_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg336_out;
SharedReg336_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg336_out;
SharedReg338_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg338_out;
SharedReg165_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg165_out;
SharedReg336_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg336_out;
   MUX_Add130_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg338_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg336_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg336_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg338_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg165_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg336_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add130_0_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_0_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Add130_1_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Add130_1_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Add130_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add130_1_impl_out,
                 X => Delay1No94_out_to_Add130_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Add130_1_impl_parent_implementedSystem_port_1_cast);

SharedReg323_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg323_out;
SharedReg325_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg325_out;
SharedReg316_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg316_out;
SharedReg323_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg323_out;
SharedReg284_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg284_out;
SharedReg15_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg15_out;
SharedReg325_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg325_out;
   MUX_Add130_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg323_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg325_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg316_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg323_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg284_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg15_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg325_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add130_1_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_1_impl_0_out,
                 Y => Delay1No94_out);

SharedReg325_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg325_out;
SharedReg337_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg337_out;
SharedReg339_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg339_out;
SharedReg325_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg325_out;
SharedReg339_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg339_out;
SharedReg31_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg31_out;
SharedReg337_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg337_out;
   MUX_Add130_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg325_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg337_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg339_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg325_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg339_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg31_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg337_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Add130_1_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_1_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Product4_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_0_impl_out,
                 X => Delay1No96_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast);

SharedReg393_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg393_out;
SharedReg396_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg67_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg67_out;
SharedReg440_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg440_out;
SharedReg39_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg39_out;
SharedReg404_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg404_out;
SharedReg38_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg38_out;
   MUX_Product4_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg393_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg67_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg440_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg39_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg404_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg38_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product4_0_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_0_out,
                 Y => Delay1No96_out);

SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg33_out;
SharedReg78_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg78_out;
SharedReg410_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg410_out;
SharedReg375_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg375_out;
SharedReg412_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg412_out;
SharedReg47_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg47_out;
SharedReg405_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg405_out;
   MUX_Product4_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg78_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg410_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg375_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg412_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg47_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg405_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product4_0_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Product4_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_1_impl_out,
                 X => Delay1No98_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg435_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg435_out;
SharedReg412_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg412_out;
SharedReg404_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg404_out;
SharedReg41_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg41_out;
SharedReg393_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg393_out;
SharedReg396_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg70_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg70_out;
   MUX_Product4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg435_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg412_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg404_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg41_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg393_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg70_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product4_1_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_0_out,
                 Y => Delay1No98_out);

SharedReg379_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg379_out;
SharedReg37_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg37_out;
SharedReg36_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg36_out;
SharedReg405_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg405_out;
SharedReg36_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg36_out;
SharedReg81_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg81_out;
SharedReg410_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg410_out;
   MUX_Product4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg379_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg37_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg36_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg405_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg36_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg81_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg410_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product4_1_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Product11_0_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Product11_0_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Product11_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_0_impl_out,
                 X => Delay1No100_out_to_Product11_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Product11_0_impl_parent_implementedSystem_port_1_cast);

SharedReg327_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg327_out;
SharedReg396_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg397_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg397_out;
SharedReg435_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg435_out;
SharedReg412_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg412_out;
SharedReg404_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg404_out;
SharedReg392_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg392_out;
   MUX_Product11_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg327_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg397_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg435_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg412_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg404_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg392_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product11_0_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_0_impl_0_out,
                 Y => Delay1No100_out);

SharedReg423_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg423_out;
SharedReg72_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg72_out;
SharedReg67_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg67_out;
SharedReg375_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg375_out;
SharedReg34_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg34_out;
SharedReg33_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg33_out;
SharedReg38_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg38_out;
   MUX_Product11_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg423_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg67_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg375_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg34_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg33_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg38_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product11_0_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_0_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Product11_1_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Product11_1_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Product11_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_1_impl_out,
                 X => Delay1No102_out_to_Product11_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Product11_1_impl_parent_implementedSystem_port_1_cast);

SharedReg147_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg147_out;
SharedReg407_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg407_out;
SharedReg395_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg395_out;
SharedReg392_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg392_out;
SharedReg332_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg332_out;
SharedReg396_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg397_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg397_out;
   MUX_Product11_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg147_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg407_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg395_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg392_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg332_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg397_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product11_1_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_1_impl_0_out,
                 Y => Delay1No102_out);

SharedReg406_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg406_out;
SharedReg106_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg106_out;
SharedReg74_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg74_out;
SharedReg41_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg41_out;
SharedReg423_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg423_out;
SharedReg75_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg75_out;
SharedReg70_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg70_out;
   MUX_Product11_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg406_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg106_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg74_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg41_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg423_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg75_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg70_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product11_1_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_1_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Product21_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_0_impl_out,
                 X => Delay1No104_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast);

SharedReg406_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg406_out;
SharedReg409_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg409_out;
SharedReg397_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg397_out;
SharedReg398_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg398_out;
SharedReg399_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg399_out;
SharedReg417_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg417_out;
SharedReg392_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg392_out;
   MUX_Product21_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg406_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg409_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg397_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg398_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg399_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg417_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg392_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product21_0_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_0_impl_0_out,
                 Y => Delay1No104_out);

SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg33_out;
SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg72_out;
SharedReg68_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg68_out;
SharedReg62_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg62_out;
SharedReg40_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg40_out;
SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg33_out;
SharedReg54_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg54_out;
   MUX_Product21_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg68_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg62_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg40_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg54_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product21_0_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_0_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Product21_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_1_impl_out,
                 X => Delay1No106_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast);

SharedReg440_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg440_out;
SharedReg42_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg42_out;
SharedReg404_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg404_out;
SharedReg392_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg392_out;
SharedReg406_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg406_out;
SharedReg409_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg409_out;
SharedReg397_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg397_out;
   MUX_Product21_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg440_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg42_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg404_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg392_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg406_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg409_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg397_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product21_1_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_1_impl_0_out,
                 Y => Delay1No106_out);

SharedReg379_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg379_out;
SharedReg412_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg412_out;
SharedReg52_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg52_out;
SharedReg57_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg57_out;
SharedReg36_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg36_out;
SharedReg75_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg75_out;
SharedReg71_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg71_out;
   MUX_Product21_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg379_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg412_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg52_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg57_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg36_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg75_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg71_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product21_1_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_1_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Subtract2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_0_impl_out,
                 X => Delay1No108_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg167_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg167_out;
SharedReg1_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg201_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg201_out;
SharedReg248_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg248_out;
SharedReg156_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg156_out;
SharedReg183_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg183_out;
SharedReg318_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg318_out;
   MUX_Subtract2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg167_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg201_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg248_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg156_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg183_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg318_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract2_0_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_0_out,
                 Y => Delay1No108_out);

SharedReg157_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg157_out;
SharedReg17_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg210_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg210_out;
SharedReg265_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg265_out;
SharedReg157_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg157_out;
SharedReg204_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg204_out;
SharedReg227_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg227_out;
   MUX_Subtract2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg157_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg210_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg265_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg157_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg204_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg227_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract2_0_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Subtract2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_1_impl_out,
                 X => Delay1No110_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg249_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg249_out;
SharedReg159_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg159_out;
SharedReg185_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg185_out;
SharedReg316_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg316_out;
SharedReg181_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg181_out;
SharedReg1_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1_out;
SharedReg208_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg208_out;
   MUX_Subtract2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg249_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg159_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg185_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg316_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg181_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg208_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract2_1_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_0_out,
                 Y => Delay1No110_out);

SharedReg267_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg267_out;
SharedReg160_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg160_out;
SharedReg207_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg207_out;
SharedReg230_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg230_out;
SharedReg160_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg160_out;
SharedReg17_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg17_out;
SharedReg225_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg225_out;
   MUX_Subtract2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg267_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg160_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg207_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg230_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg160_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg17_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg225_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract2_1_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Product5_0_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Product5_0_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Product5_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_0_impl_out,
                 X => Delay1No112_out_to_Product5_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Product5_0_impl_parent_implementedSystem_port_1_cast);

SharedReg393_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg393_out;
SharedReg78_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg78_out;
SharedReg410_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg410_out;
SharedReg411_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg411_out;
SharedReg399_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg399_out;
SharedReg402_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg402_out;
SharedReg405_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg405_out;
   MUX_Product5_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg393_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg78_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg410_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg411_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg399_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg402_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg405_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product5_0_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_0_impl_0_out,
                 Y => Delay1No112_out);

SharedReg45_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg45_out;
SharedReg409_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg409_out;
SharedReg68_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg68_out;
SharedReg62_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg62_out;
SharedReg48_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg48_out;
SharedReg44_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg44_out;
SharedReg44_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg44_out;
   MUX_Product5_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg45_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg409_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg68_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg62_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg48_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg44_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg44_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product5_0_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_0_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Product5_1_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Product5_1_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Product5_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_1_impl_out,
                 X => Delay1No114_out_to_Product5_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Product5_1_impl_parent_implementedSystem_port_1_cast);

SharedReg398_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg398_out;
SharedReg399_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg399_out;
SharedReg417_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg417_out;
SharedReg405_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg405_out;
SharedReg393_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg393_out;
SharedReg81_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg81_out;
SharedReg410_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg410_out;
   MUX_Product5_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg398_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg399_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg417_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg405_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg393_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg81_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg410_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product5_1_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_1_impl_0_out,
                 Y => Delay1No114_out);

SharedReg65_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg65_out;
SharedReg43_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg43_out;
SharedReg36_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg36_out;
SharedReg49_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg49_out;
SharedReg50_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg50_out;
SharedReg409_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg409_out;
SharedReg71_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg71_out;
   MUX_Product5_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg65_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg43_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg36_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg49_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg50_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg409_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg71_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product5_1_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_1_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Product32_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_0_impl_out,
                 X => Delay1No116_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast);

SharedReg422_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg422_out;
SharedReg396_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg397_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg397_out;
SharedReg411_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg411_out;
SharedReg412_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg412_out;
SharedReg402_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg402_out;
SharedReg54_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg54_out;
   MUX_Product32_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg422_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg397_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg411_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg412_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg402_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg54_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product32_0_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_0_out,
                 Y => Delay1No116_out);

SharedReg291_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg291_out;
SharedReg55_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg55_out;
SharedReg342_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg342_out;
SharedReg44_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg44_out;
SharedReg40_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg40_out;
SharedReg54_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg54_out;
SharedReg405_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg405_out;
   MUX_Product32_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg291_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg55_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg342_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg44_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg40_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg54_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg405_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product32_0_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Product32_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_1_impl_out,
                 X => Delay1No118_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast);

SharedReg411_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg411_out;
SharedReg399_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg399_out;
SharedReg402_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg402_out;
SharedReg57_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg57_out;
SharedReg422_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg422_out;
SharedReg396_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg397_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg397_out;
   MUX_Product32_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg411_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg399_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg402_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg57_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg422_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg397_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product32_1_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_0_out,
                 Y => Delay1No118_out);

SharedReg65_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg65_out;
SharedReg53_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg53_out;
SharedReg49_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg49_out;
SharedReg405_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg405_out;
SharedReg297_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg297_out;
SharedReg58_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg58_out;
SharedReg347_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg347_out;
   MUX_Product32_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg65_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg53_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg49_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg405_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg297_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg58_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg347_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product32_1_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Subtract3_0_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Subtract3_0_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Subtract3_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_0_impl_out,
                 X => Delay1No120_out_to_Subtract3_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Subtract3_0_impl_parent_implementedSystem_port_1_cast);

SharedReg221_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg221_out;
SharedReg2_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg2_out;
SharedReg222_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg222_out;
SharedReg228_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg228_out;
SharedReg179_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg179_out;
SharedReg227_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg227_out;
Delay5No30_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_7_cast <= Delay5No30_out;
   MUX_Subtract3_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg221_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg222_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg228_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg179_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg227_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay5No30_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract3_0_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_0_impl_0_out,
                 Y => Delay1No120_out);

SharedReg201_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg201_out;
SharedReg18_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
Delay4No12_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_3_cast <= Delay4No12_out;
SharedReg158_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg158_out;
SharedReg184_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg184_out;
SharedReg248_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg248_out;
Delay6No6_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_7_cast <= Delay6No6_out;
   MUX_Subtract3_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg201_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay4No12_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg158_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg184_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg248_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay6No6_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract3_0_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_0_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Subtract3_1_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Subtract3_1_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Subtract3_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_1_impl_out,
                 X => Delay1No122_out_to_Subtract3_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Subtract3_1_impl_parent_implementedSystem_port_1_cast);

SharedReg243_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg243_out;
SharedReg181_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg181_out;
SharedReg230_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg230_out;
Delay5No31_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_4_cast <= Delay5No31_out;
SharedReg230_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg230_out;
SharedReg2_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg2_out;
SharedReg231_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg231_out;
   MUX_Subtract3_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg243_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg181_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg230_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay5No31_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg230_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg2_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg231_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract3_1_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_1_impl_0_out,
                 Y => Delay1No122_out);

SharedReg170_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg170_out;
SharedReg186_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg186_out;
SharedReg249_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg249_out;
Delay6No7_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_4_cast <= Delay6No7_out;
SharedReg203_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg203_out;
SharedReg18_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg18_out;
Delay4No13_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_7_cast <= Delay4No13_out;
   MUX_Subtract3_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg170_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg186_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg249_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay6No7_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg203_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg18_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay4No13_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract3_1_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_1_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Product6_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_0_impl_out,
                 X => Delay1No124_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast);

SharedReg422_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg422_out;
SharedReg396_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg342_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg342_out;
SharedReg411_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg411_out;
SharedReg48_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg48_out;
SharedReg415_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg415_out;
SharedReg418_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg418_out;
   MUX_Product6_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg422_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg342_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg411_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg48_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg415_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg418_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product6_0_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_0_impl_0_out,
                 Y => Delay1No124_out);

SharedReg327_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg327_out;
SharedReg61_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg61_out;
SharedReg410_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg410_out;
SharedReg360_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg360_out;
SharedReg412_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg412_out;
SharedReg44_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg44_out;
SharedReg254_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg254_out;
   MUX_Product6_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg327_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg61_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg410_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg360_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg412_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg44_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg254_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product6_0_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_0_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Product6_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_1_impl_out,
                 X => Delay1No126_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast);

SharedReg411_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg411_out;
SharedReg412_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg412_out;
SharedReg402_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg402_out;
SharedReg418_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg418_out;
SharedReg422_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg422_out;
SharedReg396_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg347_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg347_out;
   MUX_Product6_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg411_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg412_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg402_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg418_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg422_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg347_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product6_1_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_1_impl_0_out,
                 Y => Delay1No126_out);

SharedReg49_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg49_out;
SharedReg43_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg43_out;
SharedReg57_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg57_out;
SharedReg258_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg258_out;
SharedReg332_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg332_out;
SharedReg64_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg64_out;
SharedReg410_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg410_out;
   MUX_Product6_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg49_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg43_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg57_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg258_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg332_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg64_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg410_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product6_1_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_1_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Product13_0_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Product13_0_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Product13_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product13_0_impl_out,
                 X => Delay1No128_out_to_Product13_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Product13_0_impl_parent_implementedSystem_port_1_cast);

SharedReg423_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg423_out;
SharedReg409_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg409_out;
SharedReg34_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg34_out;
SharedReg401_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg401_out;
SharedReg399_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg399_out;
SharedReg54_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg54_out;
SharedReg418_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg418_out;
   MUX_Product13_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg423_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg409_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg34_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg401_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg399_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg54_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg418_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product13_0_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_0_impl_0_out,
                 Y => Delay1No128_out);

SharedReg291_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg291_out;
SharedReg55_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg55_out;
SharedReg410_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg410_out;
SharedReg54_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg54_out;
SharedReg45_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg45_out;
SharedReg415_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg415_out;
SharedReg269_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg269_out;
   MUX_Product13_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg291_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg55_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg410_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg54_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg45_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg415_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg269_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product13_0_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_0_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Product13_1_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Product13_1_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Product13_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product13_1_impl_out,
                 X => Delay1No130_out_to_Product13_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Product13_1_impl_parent_implementedSystem_port_1_cast);

SharedReg411_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg411_out;
SharedReg53_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg53_out;
SharedReg415_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg415_out;
SharedReg418_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg418_out;
SharedReg423_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg423_out;
SharedReg409_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg409_out;
SharedReg37_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg37_out;
   MUX_Product13_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg411_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg53_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg415_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg418_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg423_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg409_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg37_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product13_1_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_1_impl_0_out,
                 Y => Delay1No130_out);

SharedReg364_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg364_out;
SharedReg412_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg412_out;
SharedReg49_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg49_out;
SharedReg273_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg273_out;
SharedReg297_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg297_out;
SharedReg58_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg58_out;
SharedReg410_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg410_out;
   MUX_Product13_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg364_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg412_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg49_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg273_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg297_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg58_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg410_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product13_1_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_1_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Product23_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_0_impl_out,
                 X => Delay1No132_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast);

SharedReg424_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg424_out;
SharedReg61_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg61_out;
SharedReg397_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg397_out;
SharedReg401_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg401_out;
SharedReg399_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg399_out;
SharedReg404_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg404_out;
SharedReg420_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg420_out;
   MUX_Product23_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg424_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg61_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg397_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg401_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg399_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg404_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg420_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product23_0_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_0_impl_0_out,
                 Y => Delay1No132_out);

SharedReg359_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg359_out;
SharedReg409_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg409_out;
SharedReg381_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg381_out;
SharedReg60_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg60_out;
SharedReg33_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg33_out;
SharedReg56_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg56_out;
SharedReg254_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg254_out;
   MUX_Product23_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg359_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg409_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg381_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg33_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg56_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg254_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product23_0_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_0_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Product23_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_1_impl_out,
                 X => Delay1No134_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast);

SharedReg401_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg401_out;
SharedReg399_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg399_out;
SharedReg57_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg57_out;
SharedReg420_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg420_out;
SharedReg424_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg424_out;
SharedReg64_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg64_out;
SharedReg397_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg397_out;
   MUX_Product23_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg401_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg399_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg57_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg420_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg424_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg64_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg397_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product23_1_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_1_impl_0_out,
                 Y => Delay1No134_out);

SharedReg57_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg57_out;
SharedReg50_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg50_out;
SharedReg415_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg415_out;
SharedReg258_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg258_out;
SharedReg363_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg363_out;
SharedReg409_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg409_out;
SharedReg384_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg384_out;
   MUX_Product23_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg57_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg50_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg415_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg258_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg363_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg409_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg384_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product23_1_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_1_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Product33_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_0_impl_out,
                 X => Delay1No136_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast);

SharedReg424_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg424_out;
SharedReg396_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg381_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg381_out;
SharedReg414_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg414_out;
SharedReg33_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg33_out;
SharedReg417_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg417_out;
SharedReg269_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg269_out;
   MUX_Product33_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg424_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg381_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg414_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg33_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg417_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg269_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product33_0_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_0_impl_0_out,
                 Y => Delay1No136_out);

SharedReg341_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg341_out;
SharedReg73_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg73_out;
SharedReg410_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg410_out;
SharedReg54_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg54_out;
SharedReg412_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg412_out;
SharedReg56_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg56_out;
SharedReg420_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg420_out;
   MUX_Product33_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg341_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg73_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg410_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg54_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg412_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg56_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg420_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product33_0_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_0_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Product33_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_1_impl_out,
                 X => Delay1No138_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast);

SharedReg401_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg401_out;
SharedReg399_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg399_out;
SharedReg404_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg404_out;
SharedReg273_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg273_out;
SharedReg424_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg424_out;
SharedReg396_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg384_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg384_out;
   MUX_Product33_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg401_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg399_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg404_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg273_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg424_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg384_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product33_1_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_1_impl_0_out,
                 Y => Delay1No138_out);

SharedReg63_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg63_out;
SharedReg36_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg36_out;
SharedReg59_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg59_out;
SharedReg420_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg420_out;
SharedReg346_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg346_out;
SharedReg76_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg76_out;
SharedReg410_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg410_out;
   MUX_Product33_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg63_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg36_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg59_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg420_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg346_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg76_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg410_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product33_1_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_1_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Subtract4_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_0_impl_out,
                 X => Delay1No140_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast);

SharedReg162_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg162_out;
SharedReg_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg168_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg168_out;
SharedReg195_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg195_out;
SharedReg183_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg183_out;
SharedReg162_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg162_out;
SharedReg167_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg167_out;
   MUX_Subtract4_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg162_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg168_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg195_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg183_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg162_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg167_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract4_0_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_0_impl_0_out,
                 Y => Delay1No140_out);

SharedReg229_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg229_out;
SharedReg16_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg196_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg196_out;
SharedReg209_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg209_out;
SharedReg162_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg162_out;
SharedReg179_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg179_out;
SharedReg222_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg222_out;
   MUX_Subtract4_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg229_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg196_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg209_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg162_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg179_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg222_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract4_0_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_0_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Subtract4_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_1_impl_out,
                 X => Delay1No142_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg197_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg197_out;
SharedReg185_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg185_out;
SharedReg165_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg165_out;
SharedReg169_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg169_out;
SharedReg159_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg159_out;
SharedReg_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg_out;
SharedReg182_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg182_out;
   MUX_Subtract4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg197_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg185_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg165_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg169_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg159_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg182_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract4_1_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_1_impl_0_out,
                 Y => Delay1No142_out);

SharedReg212_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg212_out;
SharedReg165_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg165_out;
SharedReg181_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg181_out;
SharedReg225_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg225_out;
SharedReg232_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg232_out;
SharedReg16_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg16_out;
SharedReg203_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg203_out;
   MUX_Subtract4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg212_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg165_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg181_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg225_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg232_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg16_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg203_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract4_1_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_1_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Product25_0_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Product25_0_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Product25_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product25_0_impl_out,
                 X => Delay1No144_out_to_Product25_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Product25_0_impl_parent_implementedSystem_port_1_cast);

SharedReg428_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg428_out;
SharedReg73_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg73_out;
SharedReg437_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg437_out;
SharedReg398_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg398_out;
SharedReg399_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg399_out;
SharedReg404_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg404_out;
SharedReg434_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg434_out;
   MUX_Product25_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg428_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg73_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg437_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg398_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg399_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg404_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg434_out_to_MUX_Product25_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product25_0_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product25_0_impl_0_out,
                 Y => Delay1No144_out);

SharedReg359_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg359_out;
SharedReg409_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg409_out;
SharedReg382_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg382_out;
SharedReg34_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg34_out;
SharedReg361_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg361_out;
SharedReg368_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg368_out;
SharedReg380_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg380_out;
   MUX_Product25_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg359_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg409_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg382_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg34_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg361_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg368_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg380_out_to_MUX_Product25_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product25_0_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product25_0_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Product25_1_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Product25_1_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Product25_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product25_1_impl_out,
                 X => Delay1No146_out_to_Product25_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Product25_1_impl_parent_implementedSystem_port_1_cast);

SharedReg414_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg414_out;
SharedReg36_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg36_out;
SharedReg417_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg417_out;
SharedReg434_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg434_out;
SharedReg428_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg428_out;
SharedReg76_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg76_out;
SharedReg437_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg437_out;
   MUX_Product25_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg414_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg36_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg417_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg434_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg428_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg76_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg437_out_to_MUX_Product25_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product25_1_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product25_1_impl_0_out,
                 Y => Delay1No146_out);

SharedReg57_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg57_out;
SharedReg412_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg412_out;
SharedReg59_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg59_out;
SharedReg383_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg383_out;
SharedReg363_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg363_out;
SharedReg409_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg409_out;
SharedReg385_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg385_out;
   MUX_Product25_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg57_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg412_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg59_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg383_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg363_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg409_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg385_out_to_MUX_Product25_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product25_1_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product25_1_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Product35_0_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Product35_0_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Product35_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product35_0_impl_out,
                 X => Delay1No148_out_to_Product35_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Product35_0_impl_parent_implementedSystem_port_1_cast);

SharedReg341_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg341_out;
SharedReg419_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg419_out;
SharedReg382_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg382_out;
SharedReg411_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg411_out;
SharedReg399_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg399_out;
SharedReg417_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg417_out;
SharedReg380_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg380_out;
   MUX_Product35_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg341_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg419_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg382_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg411_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg399_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg417_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg380_out_to_MUX_Product35_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product35_0_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product35_0_impl_0_out,
                 Y => Delay1No148_out);

SharedReg428_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg428_out;
SharedReg351_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg351_out;
SharedReg442_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg442_out;
SharedReg34_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg34_out;
SharedReg34_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg34_out;
SharedReg368_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg368_out;
SharedReg439_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg439_out;
   MUX_Product35_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg428_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg351_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg442_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg34_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg34_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg368_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg439_out_to_MUX_Product35_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product35_0_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product35_0_impl_1_out,
                 Y => Delay1No149_out);

Delay1No150_out_to_Product35_1_impl_parent_implementedSystem_port_0_cast <= Delay1No150_out;
Delay1No151_out_to_Product35_1_impl_parent_implementedSystem_port_1_cast <= Delay1No151_out;
   Product35_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product35_1_impl_out,
                 X => Delay1No150_out_to_Product35_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No151_out_to_Product35_1_impl_parent_implementedSystem_port_1_cast);

SharedReg398_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg398_out;
SharedReg399_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg399_out;
SharedReg404_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg404_out;
SharedReg383_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg383_out;
SharedReg346_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg346_out;
SharedReg419_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg419_out;
SharedReg385_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg385_out;
   MUX_Product35_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg398_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg399_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg404_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg383_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg346_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg419_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg385_out_to_MUX_Product35_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product35_1_impl_0_out);

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product35_1_impl_0_out,
                 Y => Delay1No150_out);

SharedReg37_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg37_out;
SharedReg365_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg365_out;
SharedReg371_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg371_out;
SharedReg439_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg439_out;
SharedReg428_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg428_out;
SharedReg355_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg355_out;
SharedReg442_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg442_out;
   MUX_Product35_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg37_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg365_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg371_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg439_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg428_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg355_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg442_out_to_MUX_Product35_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product35_1_impl_1_out);

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product35_1_impl_1_out,
                 Y => Delay1No151_out);

Delay1No152_out_to_Subtract6_0_impl_parent_implementedSystem_port_0_cast <= Delay1No152_out;
Delay1No153_out_to_Subtract6_0_impl_parent_implementedSystem_port_1_cast <= Delay1No153_out;
   Subtract6_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract6_0_impl_out,
                 X => Delay1No152_out_to_Subtract6_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No153_out_to_Subtract6_0_impl_parent_implementedSystem_port_1_cast);

SharedReg239_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg239_out;
SharedReg3_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg286_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg286_out;
Delay3No66_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_4_cast <= Delay3No66_out;
SharedReg204_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg204_out;
SharedReg262_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg262_out;
SharedReg223_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg223_out;
   MUX_Subtract6_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg239_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg286_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay3No66_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg204_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg262_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg223_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract6_0_impl_0_out);

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_0_impl_0_out,
                 Y => Delay1No152_out);

Delay3No86_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_1_cast <= Delay3No86_out;
SharedReg19_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg312_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg312_out;
Delay5No28_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_4_cast <= Delay5No28_out;
SharedReg227_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg227_out;
SharedReg285_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg285_out;
Delay6No10_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_7_cast <= Delay6No10_out;
   MUX_Subtract6_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No86_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg312_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay5No28_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg227_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg285_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay6No10_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract6_0_impl_1_out);

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_0_impl_1_out,
                 Y => Delay1No153_out);

Delay1No154_out_to_Subtract6_1_impl_parent_implementedSystem_port_0_cast <= Delay1No154_out;
Delay1No155_out_to_Subtract6_1_impl_parent_implementedSystem_port_1_cast <= Delay1No155_out;
   Subtract6_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract6_1_impl_out,
                 X => Delay1No154_out_to_Subtract6_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No155_out_to_Subtract6_1_impl_parent_implementedSystem_port_1_cast);

Delay3No67_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_1_cast <= Delay3No67_out;
SharedReg207_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg207_out;
SharedReg264_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg264_out;
SharedReg232_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg232_out;
SharedReg246_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg246_out;
SharedReg3_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg3_out;
SharedReg305_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg305_out;
   MUX_Subtract6_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No67_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg207_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg264_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg232_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg246_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg3_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg305_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract6_1_impl_0_out);

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_1_impl_0_out,
                 Y => Delay1No154_out);

Delay5No29_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_1_cast <= Delay5No29_out;
SharedReg230_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg230_out;
SharedReg288_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg288_out;
Delay6No11_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_4_cast <= Delay6No11_out;
Delay3No87_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_5_cast <= Delay3No87_out;
SharedReg19_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg19_out;
SharedReg316_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg316_out;
   MUX_Subtract6_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No29_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg230_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg288_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay6No11_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay3No87_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg19_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg316_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract6_1_impl_1_out);

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_1_impl_1_out,
                 Y => Delay1No155_out);

Delay1No156_out_to_Product9_0_impl_parent_implementedSystem_port_0_cast <= Delay1No156_out;
Delay1No157_out_to_Product9_0_impl_parent_implementedSystem_port_1_cast <= Delay1No157_out;
   Product9_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product9_0_impl_out,
                 X => Delay1No156_out_to_Product9_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No157_out_to_Product9_0_impl_parent_implementedSystem_port_1_cast);

SharedReg432_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg432_out;
SharedReg419_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg419_out;
SharedReg400_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg400_out;
SharedReg438_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg438_out;
SharedReg399_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg399_out;
SharedReg402_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg402_out;
SharedReg444_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg444_out;
   MUX_Product9_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg432_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg419_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg400_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg438_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg399_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg402_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg444_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product9_0_impl_0_out);

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_0_impl_0_out,
                 Y => Delay1No156_out);

SharedReg351_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg351_out;
SharedReg367_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg367_out;
SharedReg66_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg66_out;
SharedReg328_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg328_out;
SharedReg39_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg39_out;
SharedReg32_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg32_out;
SharedReg390_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg390_out;
   MUX_Product9_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg351_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg367_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg66_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg328_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg39_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg32_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg390_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product9_0_impl_1_out);

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_0_impl_1_out,
                 Y => Delay1No157_out);

Delay1No158_out_to_Product9_1_impl_parent_implementedSystem_port_0_cast <= Delay1No158_out;
Delay1No159_out_to_Product9_1_impl_parent_implementedSystem_port_1_cast <= Delay1No159_out;
   Product9_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product9_1_impl_out,
                 X => Delay1No158_out_to_Product9_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No159_out_to_Product9_1_impl_parent_implementedSystem_port_1_cast);

SharedReg411_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg411_out;
SharedReg399_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg399_out;
SharedReg417_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg417_out;
SharedReg444_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg444_out;
SharedReg432_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg432_out;
SharedReg419_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg419_out;
SharedReg400_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg400_out;
   MUX_Product9_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg411_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg399_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg417_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg444_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg432_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg419_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg400_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product9_1_impl_0_out);

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_1_impl_0_out,
                 Y => Delay1No158_out);

SharedReg37_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg37_out;
SharedReg37_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg37_out;
SharedReg371_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg371_out;
SharedReg391_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg391_out;
SharedReg355_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg355_out;
SharedReg370_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg370_out;
SharedReg69_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg69_out;
   MUX_Product9_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg37_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg37_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg371_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg391_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg355_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg370_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg69_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product9_1_impl_1_out);

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_1_impl_1_out,
                 Y => Delay1No159_out);

Delay1No160_out_to_Product16_0_impl_parent_implementedSystem_port_0_cast <= Delay1No160_out;
Delay1No161_out_to_Product16_0_impl_parent_implementedSystem_port_1_cast <= Delay1No161_out;
   Product16_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product16_0_impl_out,
                 X => Delay1No160_out_to_Product16_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No161_out_to_Product16_0_impl_parent_implementedSystem_port_1_cast);

SharedReg432_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg432_out;
SharedReg421_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg421_out;
SharedReg400_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg400_out;
SharedReg443_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg443_out;
SharedReg399_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg399_out;
SharedReg402_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg402_out;
SharedReg390_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg390_out;
   MUX_Product16_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg432_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg421_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg400_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg443_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg399_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg402_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg390_out_to_MUX_Product16_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product16_0_impl_0_out);

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product16_0_impl_0_out,
                 Y => Delay1No160_out);

SharedReg367_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg367_out;
SharedReg351_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg351_out;
SharedReg72_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg72_out;
SharedReg328_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg328_out;
SharedReg374_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg374_out;
SharedReg38_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg38_out;
SharedReg446_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg446_out;
   MUX_Product16_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg367_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg351_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg72_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg328_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg374_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg38_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg446_out_to_MUX_Product16_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product16_0_impl_1_out);

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product16_0_impl_1_out,
                 Y => Delay1No161_out);

Delay1No162_out_to_Product16_1_impl_parent_implementedSystem_port_0_cast <= Delay1No162_out;
Delay1No163_out_to_Product16_1_impl_parent_implementedSystem_port_1_cast <= Delay1No163_out;
   Product16_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product16_1_impl_out,
                 X => Delay1No162_out_to_Product16_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No163_out_to_Product16_1_impl_parent_implementedSystem_port_1_cast);

SharedReg438_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg438_out;
SharedReg399_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg399_out;
SharedReg402_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg402_out;
SharedReg391_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg391_out;
SharedReg432_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg432_out;
SharedReg421_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg421_out;
SharedReg400_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg400_out;
   MUX_Product16_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg438_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg399_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg402_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg391_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg432_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg421_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg400_out_to_MUX_Product16_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product16_1_impl_0_out);

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product16_1_impl_0_out,
                 Y => Delay1No162_out);

SharedReg333_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg333_out;
SharedReg42_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg42_out;
SharedReg35_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg35_out;
SharedReg446_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg446_out;
SharedReg370_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg370_out;
SharedReg355_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg355_out;
SharedReg75_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg75_out;
   MUX_Product16_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg333_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg42_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg35_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg446_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg370_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg355_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg75_out_to_MUX_Product16_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product16_1_impl_1_out);

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product16_1_impl_1_out,
                 Y => Delay1No163_out);

Delay1No164_out_to_Product26_0_impl_parent_implementedSystem_port_0_cast <= Delay1No164_out;
Delay1No165_out_to_Product26_0_impl_parent_implementedSystem_port_1_cast <= Delay1No165_out;
   Product26_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_0_impl_out,
                 X => Delay1No164_out_to_Product26_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No165_out_to_Product26_0_impl_parent_implementedSystem_port_1_cast);

SharedReg433_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg433_out;
SharedReg367_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg367_out;
SharedReg413_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg413_out;
SharedReg60_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg60_out;
SharedReg412_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg412_out;
SharedReg415_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg415_out;
SharedReg392_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg392_out;
   MUX_Product26_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg433_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg367_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg413_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg412_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg415_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg392_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product26_0_impl_0_out);

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_0_impl_0_out,
                 Y => Delay1No164_out);

SharedReg351_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg351_out;
SharedReg421_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg421_out;
SharedReg66_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg66_out;
SharedReg414_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg414_out;
SharedReg374_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg374_out;
SharedReg32_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg32_out;
SharedReg60_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg60_out;
   MUX_Product26_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg351_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg421_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg66_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg414_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg374_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg32_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg60_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product26_0_impl_1_out);

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_0_impl_1_out,
                 Y => Delay1No165_out);

Delay1No166_out_to_Product26_1_impl_parent_implementedSystem_port_0_cast <= Delay1No166_out;
Delay1No167_out_to_Product26_1_impl_parent_implementedSystem_port_1_cast <= Delay1No167_out;
   Product26_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_1_impl_out,
                 X => Delay1No166_out_to_Product26_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No167_out_to_Product26_1_impl_parent_implementedSystem_port_1_cast);

SharedReg443_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg443_out;
SharedReg399_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg399_out;
SharedReg402_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg402_out;
SharedReg392_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg392_out;
SharedReg433_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg433_out;
SharedReg370_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg370_out;
SharedReg413_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg413_out;
   MUX_Product26_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg443_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg399_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg402_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg392_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg433_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg370_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg413_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product26_1_impl_0_out);

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_1_impl_0_out,
                 Y => Delay1No166_out);

SharedReg333_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg333_out;
SharedReg378_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg378_out;
SharedReg41_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg41_out;
SharedReg63_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg63_out;
SharedReg355_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg355_out;
SharedReg421_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg421_out;
SharedReg69_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg69_out;
   MUX_Product26_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg333_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg378_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg41_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg63_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg355_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg421_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg69_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product26_1_impl_1_out);

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_1_impl_1_out,
                 Y => Delay1No167_out);

Delay1No168_out_to_Product36_0_impl_parent_implementedSystem_port_0_cast <= Delay1No168_out;
Delay1No169_out_to_Product36_0_impl_parent_implementedSystem_port_1_cast <= Delay1No169_out;
   Product36_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product36_0_impl_out,
                 X => Delay1No168_out_to_Product36_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No169_out_to_Product36_0_impl_parent_implementedSystem_port_1_cast);

SharedReg367_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg367_out;
SharedReg396_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg72_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg72_out;
SharedReg401_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg401_out;
SharedReg425_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg425_out;
SharedReg38_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg38_out;
SharedReg392_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg392_out;
   MUX_Product36_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg367_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg72_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg401_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg425_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg38_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg392_out_to_MUX_Product36_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product36_0_impl_0_out);

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product36_0_impl_0_out,
                 Y => Delay1No168_out);

SharedReg433_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg433_out;
SharedReg33_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg33_out;
SharedReg413_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg413_out;
SharedReg66_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg66_out;
SharedReg352_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg352_out;
SharedReg415_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg415_out;
SharedReg66_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg66_out;
   MUX_Product36_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg433_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg33_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg413_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg66_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg352_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg415_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg66_out_to_MUX_Product36_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product36_0_impl_1_out);

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product36_0_impl_1_out,
                 Y => Delay1No169_out);

Delay1No170_out_to_Product36_1_impl_parent_implementedSystem_port_0_cast <= Delay1No170_out;
Delay1No171_out_to_Product36_1_impl_parent_implementedSystem_port_1_cast <= Delay1No171_out;
   Product36_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product36_1_impl_out,
                 X => Delay1No170_out_to_Product36_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No171_out_to_Product36_1_impl_parent_implementedSystem_port_1_cast);

SharedReg63_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg63_out;
SharedReg412_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg412_out;
SharedReg415_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg415_out;
SharedReg392_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg392_out;
SharedReg370_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg370_out;
SharedReg396_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg75_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg75_out;
   MUX_Product36_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg63_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg412_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg415_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg392_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg370_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg75_out_to_MUX_Product36_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product36_1_impl_0_out);

   Delay1No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product36_1_impl_0_out,
                 Y => Delay1No170_out);

SharedReg414_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg414_out;
SharedReg378_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg378_out;
SharedReg35_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg35_out;
SharedReg69_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg69_out;
SharedReg433_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg433_out;
SharedReg36_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg36_out;
SharedReg413_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg413_out;
   MUX_Product36_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg414_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg378_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg35_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg69_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg433_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg36_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg413_out_to_MUX_Product36_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product36_1_impl_1_out);

   Delay1No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product36_1_impl_1_out,
                 Y => Delay1No171_out);

Delay1No172_out_to_Subtract7_0_impl_parent_implementedSystem_port_0_cast <= Delay1No172_out;
Delay1No173_out_to_Subtract7_0_impl_parent_implementedSystem_port_1_cast <= Delay1No173_out;
   Subtract7_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract7_0_impl_out,
                 X => Delay1No172_out_to_Subtract7_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No173_out_to_Subtract7_0_impl_parent_implementedSystem_port_1_cast);

SharedReg200_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg200_out;
SharedReg4_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg4_out;
SharedReg239_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg239_out;
SharedReg180_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg180_out;
SharedReg239_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg239_out;
SharedReg278_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg278_out;
SharedReg239_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg239_out;
   MUX_Subtract7_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg200_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg4_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg239_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg180_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg239_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg278_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg239_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract7_0_impl_0_out);

   Delay1No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_0_impl_0_out,
                 Y => Delay1No172_out);

SharedReg248_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg248_out;
SharedReg20_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg250_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg250_out;
SharedReg201_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg201_out;
SharedReg250_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg250_out;
SharedReg311_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg311_out;
SharedReg250_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg250_out;
   MUX_Subtract7_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg248_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg250_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg201_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg250_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg311_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg250_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract7_0_impl_1_out);

   Delay1No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_0_impl_1_out,
                 Y => Delay1No173_out);

Delay1No174_out_to_Subtract7_1_impl_parent_implementedSystem_port_0_cast <= Delay1No174_out;
Delay1No175_out_to_Subtract7_1_impl_parent_implementedSystem_port_1_cast <= Delay1No175_out;
   Subtract7_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract7_1_impl_out,
                 X => Delay1No174_out_to_Subtract7_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No175_out_to_Subtract7_1_impl_parent_implementedSystem_port_1_cast);

SharedReg186_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg186_out;
SharedReg241_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg241_out;
SharedReg282_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg282_out;
SharedReg241_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg241_out;
SharedReg207_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg207_out;
SharedReg4_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg4_out;
SharedReg246_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg246_out;
   MUX_Subtract7_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg186_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg241_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg282_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg241_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg207_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg4_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg246_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract7_1_impl_0_out);

   Delay1No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_1_impl_0_out,
                 Y => Delay1No174_out);

SharedReg208_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg208_out;
SharedReg252_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg252_out;
SharedReg313_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg313_out;
SharedReg252_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg252_out;
SharedReg252_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg252_out;
SharedReg20_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg20_out;
SharedReg264_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg264_out;
   MUX_Subtract7_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg208_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg252_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg313_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg252_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg252_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg20_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg264_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract7_1_impl_1_out);

   Delay1No175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_1_impl_1_out,
                 Y => Delay1No175_out);

Delay1No176_out_to_Product18_0_impl_parent_implementedSystem_port_0_cast <= Delay1No176_out;
Delay1No177_out_to_Product18_0_impl_parent_implementedSystem_port_1_cast <= Delay1No177_out;
   Product18_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_0_impl_out,
                 X => Delay1No176_out_to_Product18_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No177_out_to_Product18_0_impl_parent_implementedSystem_port_1_cast);

SharedReg445_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg445_out;
SharedReg419_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg419_out;
SharedReg426_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg426_out;
SharedReg401_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg401_out;
SharedReg425_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg425_out;
SharedReg404_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg404_out;
SharedReg405_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg405_out;
   MUX_Product18_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg445_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg419_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg426_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg401_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg425_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg404_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg405_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product18_0_impl_0_out);

   Delay1No176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_0_impl_0_out,
                 Y => Delay1No176_out);

SharedReg387_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg387_out;
SharedReg386_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg386_out;
SharedReg372_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg372_out;
SharedReg72_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg72_out;
SharedReg341_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg341_out;
SharedReg373_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg373_out;
SharedReg60_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg60_out;
   MUX_Product18_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg387_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg386_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg372_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg72_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg341_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg373_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg60_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product18_0_impl_1_out);

   Delay1No177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_0_impl_1_out,
                 Y => Delay1No177_out);

Delay1No178_out_to_Product18_1_impl_parent_implementedSystem_port_0_cast <= Delay1No178_out;
Delay1No179_out_to_Product18_1_impl_parent_implementedSystem_port_1_cast <= Delay1No179_out;
   Product18_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_1_impl_out,
                 X => Delay1No178_out_to_Product18_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No179_out_to_Product18_1_impl_parent_implementedSystem_port_1_cast);

SharedReg401_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg401_out;
SharedReg425_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg425_out;
SharedReg41_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg41_out;
SharedReg405_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg405_out;
SharedReg445_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg445_out;
SharedReg419_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg419_out;
SharedReg426_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg426_out;
   MUX_Product18_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg401_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg425_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg41_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg405_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg445_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg419_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg426_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product18_1_impl_0_out);

   Delay1No178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_1_impl_0_out,
                 Y => Delay1No178_out);

SharedReg69_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg69_out;
SharedReg356_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg356_out;
SharedReg415_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg415_out;
SharedReg63_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg63_out;
SharedReg389_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg389_out;
SharedReg388_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg388_out;
SharedReg376_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg376_out;
   MUX_Product18_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg356_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg415_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg63_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg389_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg388_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg376_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product18_1_impl_1_out);

   Delay1No179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_1_impl_1_out,
                 Y => Delay1No179_out);

Delay1No180_out_to_Product28_0_impl_parent_implementedSystem_port_0_cast <= Delay1No180_out;
Delay1No181_out_to_Product28_0_impl_parent_implementedSystem_port_1_cast <= Delay1No181_out;
   Product28_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_0_impl_out,
                 X => Delay1No180_out_to_Product28_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No181_out_to_Product28_0_impl_parent_implementedSystem_port_1_cast);

SharedReg447_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg447_out;
SharedReg419_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg419_out;
SharedReg426_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg426_out;
SharedReg414_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg414_out;
SharedReg429_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg429_out;
SharedReg404_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg404_out;
SharedReg66_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg66_out;
   MUX_Product28_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg447_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg419_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg426_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg414_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg429_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg404_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg66_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product28_0_impl_0_out);

   Delay1No180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_0_impl_0_out,
                 Y => Delay1No180_out);

SharedReg387_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg387_out;
SharedReg390_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg390_out;
SharedReg380_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg380_out;
SharedReg66_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg66_out;
SharedReg352_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg352_out;
SharedReg361_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg361_out;
SharedReg405_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg405_out;
   MUX_Product28_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg387_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg390_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg380_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg66_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg352_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg361_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg405_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product28_0_impl_1_out);

   Delay1No181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_0_impl_1_out,
                 Y => Delay1No181_out);

Delay1No182_out_to_Product28_1_impl_parent_implementedSystem_port_0_cast <= Delay1No182_out;
Delay1No183_out_to_Product28_1_impl_parent_implementedSystem_port_1_cast <= Delay1No183_out;
   Product28_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_1_impl_out,
                 X => Delay1No182_out_to_Product28_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No183_out_to_Product28_1_impl_parent_implementedSystem_port_1_cast);

SharedReg401_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg401_out;
SharedReg425_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg425_out;
SharedReg404_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg404_out;
SharedReg69_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg69_out;
SharedReg447_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg447_out;
SharedReg419_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg419_out;
SharedReg426_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg426_out;
   MUX_Product28_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg401_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg425_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg404_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg69_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg447_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg419_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg426_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product28_1_impl_0_out);

   Delay1No182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_1_impl_0_out,
                 Y => Delay1No182_out);

SharedReg75_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg75_out;
SharedReg346_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg346_out;
SharedReg377_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg377_out;
SharedReg405_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg405_out;
SharedReg389_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg389_out;
SharedReg391_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg391_out;
SharedReg383_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg383_out;
   MUX_Product28_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg75_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg346_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg377_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg405_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg389_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg391_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg383_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product28_1_impl_1_out);

   Delay1No183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_1_impl_1_out,
                 Y => Delay1No183_out);

Delay1No184_out_to_Subtract9_0_impl_parent_implementedSystem_port_0_cast <= Delay1No184_out;
Delay1No185_out_to_Subtract9_0_impl_parent_implementedSystem_port_1_cast <= Delay1No185_out;
   Subtract9_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_0_impl_out,
                 X => Delay1No184_out_to_Subtract9_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No185_out_to_Subtract9_0_impl_parent_implementedSystem_port_1_cast);

SharedReg250_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg250_out;
SharedReg5_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg302_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg302_out;
SharedReg302_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg302_out;
SharedReg262_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg262_out;
SharedReg324_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg324_out;
Delay5No42_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_7_cast <= Delay5No42_out;
   MUX_Subtract9_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg250_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg302_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg302_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg262_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg324_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay5No42_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract9_0_impl_0_out);

   Delay1No184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_0_impl_0_out,
                 Y => Delay1No184_out);

SharedReg277_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg277_out;
SharedReg21_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg21_out;
SharedReg317_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg317_out;
SharedReg245_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg245_out;
SharedReg312_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg312_out;
Delay5No48_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_7_cast <= Delay5No48_out;
   MUX_Subtract9_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg277_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg21_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg317_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg317_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg245_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg312_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay5No48_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract9_0_impl_1_out);

   Delay1No185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_0_impl_1_out,
                 Y => Delay1No185_out);

Delay1No186_out_to_Subtract9_1_impl_parent_implementedSystem_port_0_cast <= Delay1No186_out;
Delay1No187_out_to_Subtract9_1_impl_parent_implementedSystem_port_1_cast <= Delay1No187_out;
   Subtract9_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_1_impl_out,
                 X => Delay1No186_out_to_Subtract9_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No187_out_to_Subtract9_1_impl_parent_implementedSystem_port_1_cast);

SharedReg304_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg304_out;
SharedReg264_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg264_out;
SharedReg323_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg323_out;
Delay5No43_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_4_cast <= Delay5No43_out;
SharedReg264_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg264_out;
SharedReg5_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg5_out;
SharedReg309_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg309_out;
   MUX_Subtract9_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg304_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg264_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg323_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay5No43_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg264_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg5_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg309_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract9_1_impl_0_out);

   Delay1No186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_1_impl_0_out,
                 Y => Delay1No186_out);

SharedReg315_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg315_out;
SharedReg247_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg247_out;
SharedReg314_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg314_out;
Delay5No49_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_4_cast <= Delay5No49_out;
SharedReg288_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg288_out;
SharedReg21_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg21_out;
SharedReg321_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg321_out;
   MUX_Subtract9_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg315_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg247_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg314_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay5No49_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg288_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg21_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg321_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract9_1_impl_1_out);

   Delay1No187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_1_impl_1_out,
                 Y => Delay1No187_out);

Delay1No188_out_to_Product221_0_impl_parent_implementedSystem_port_0_cast <= Delay1No188_out;
Delay1No189_out_to_Product221_0_impl_parent_implementedSystem_port_1_cast <= Delay1No189_out;
   Product221_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_0_impl_out,
                 X => Delay1No188_out_to_Product221_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No189_out_to_Product221_0_impl_parent_implementedSystem_port_1_cast);

SharedReg393_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg393_out;
SharedReg421_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg421_out;
SharedReg430_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg430_out;
SharedReg72_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg72_out;
SharedReg341_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg341_out;
SharedReg417_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg417_out;
SharedReg392_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg392_out;
   MUX_Product221_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg393_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg421_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg430_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg72_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg341_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg417_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg392_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product221_0_impl_0_out);

   Delay1No188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_0_impl_0_out,
                 Y => Delay1No188_out);

SharedReg79_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg79_out;
SharedReg386_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg386_out;
SharedReg372_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg372_out;
SharedReg414_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg414_out;
SharedReg429_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg429_out;
SharedReg373_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg373_out;
SharedReg124_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg124_out;
   MUX_Product221_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg79_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg386_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg372_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg414_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg429_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg373_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg124_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product221_0_impl_1_out);

   Delay1No189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_0_impl_1_out,
                 Y => Delay1No189_out);

Delay1No190_out_to_Product221_1_impl_parent_implementedSystem_port_0_cast <= Delay1No190_out;
Delay1No191_out_to_Product221_1_impl_parent_implementedSystem_port_1_cast <= Delay1No191_out;
   Product221_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_1_impl_out,
                 X => Delay1No190_out_to_Product221_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No191_out_to_Product221_1_impl_parent_implementedSystem_port_1_cast);

SharedReg414_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg414_out;
SharedReg429_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg429_out;
SharedReg404_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg404_out;
SharedReg392_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg392_out;
SharedReg393_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg393_out;
SharedReg421_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg421_out;
SharedReg430_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg430_out;
   MUX_Product221_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg414_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg429_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg404_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg392_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg393_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg421_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg430_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product221_1_impl_0_out);

   Delay1No190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_1_impl_0_out,
                 Y => Delay1No190_out);

SharedReg69_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg69_out;
SharedReg356_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg356_out;
SharedReg365_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg365_out;
SharedReg130_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg130_out;
SharedReg82_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg82_out;
SharedReg388_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg388_out;
SharedReg376_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg376_out;
   MUX_Product221_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg356_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg365_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg130_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg82_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg388_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg376_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product221_1_impl_1_out);

   Delay1No191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_1_impl_1_out,
                 Y => Delay1No191_out);

Delay1No192_out_to_Product321_0_impl_parent_implementedSystem_port_0_cast <= Delay1No192_out;
Delay1No193_out_to_Product321_0_impl_parent_implementedSystem_port_1_cast <= Delay1No193_out;
   Product321_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_0_impl_out,
                 X => Delay1No192_out_to_Product321_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No193_out_to_Product321_0_impl_parent_implementedSystem_port_1_cast);

SharedReg393_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg393_out;
SharedReg390_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg390_out;
SharedReg380_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg380_out;
SharedReg427_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg427_out;
SharedReg425_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg425_out;
SharedReg361_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg361_out;
SharedReg124_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg124_out;
   MUX_Product321_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg393_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg390_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg380_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg427_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg425_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg361_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg124_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product321_0_impl_0_out);

   Delay1No192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_0_impl_0_out,
                 Y => Delay1No192_out);

SharedReg85_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg85_out;
SharedReg421_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg421_out;
SharedReg430_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg430_out;
SharedReg386_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg386_out;
SharedReg351_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg351_out;
SharedReg417_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg417_out;
SharedReg405_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg405_out;
   MUX_Product321_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg85_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg421_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg430_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg386_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg351_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg417_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg405_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product321_0_impl_1_out);

   Delay1No193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_0_impl_1_out,
                 Y => Delay1No193_out);

Delay1No194_out_to_Product321_1_impl_parent_implementedSystem_port_0_cast <= Delay1No194_out;
Delay1No195_out_to_Product321_1_impl_parent_implementedSystem_port_1_cast <= Delay1No195_out;
   Product321_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_1_impl_out,
                 X => Delay1No194_out_to_Product321_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No195_out_to_Product321_1_impl_parent_implementedSystem_port_1_cast);

SharedReg75_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg75_out;
SharedReg346_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg346_out;
SharedReg417_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg417_out;
SharedReg130_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg130_out;
SharedReg393_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg393_out;
SharedReg391_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg391_out;
SharedReg383_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg383_out;
   MUX_Product321_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg75_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg346_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg417_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg130_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg393_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg391_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg383_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product321_1_impl_0_out);

   Delay1No194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_1_impl_0_out,
                 Y => Delay1No194_out);

SharedReg414_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg414_out;
SharedReg429_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg429_out;
SharedReg377_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg377_out;
SharedReg405_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg405_out;
SharedReg88_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg88_out;
SharedReg421_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg421_out;
SharedReg430_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg430_out;
   MUX_Product321_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg414_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg429_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg377_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg405_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg88_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg421_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg430_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product321_1_impl_1_out);

   Delay1No195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_1_impl_1_out,
                 Y => Delay1No195_out);

Delay1No196_out_to_Subtract23_0_impl_parent_implementedSystem_port_0_cast <= Delay1No196_out;
Delay1No197_out_to_Subtract23_0_impl_parent_implementedSystem_port_1_cast <= Delay1No197_out;
   Subtract23_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract23_0_impl_out,
                 X => Delay1No196_out_to_Subtract23_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No197_out_to_Subtract23_0_impl_parent_implementedSystem_port_1_cast);

SharedReg285_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg285_out;
SharedReg6_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg6_out;
SharedReg319_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg319_out;
SharedReg319_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg319_out;
Delay4No22_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_5_cast <= Delay4No22_out;
SharedReg126_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg126_out;
SharedReg262_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg262_out;
   MUX_Subtract23_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg285_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg6_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg319_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg319_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay4No22_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg126_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg262_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract23_0_impl_0_out);

   Delay1No196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_0_impl_0_out,
                 Y => Delay1No196_out);

SharedReg311_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg311_out;
SharedReg22_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg22_out;
SharedReg338_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg338_out;
SharedReg279_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg279_out;
SharedReg118_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg118_out;
SharedReg285_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg285_out;
   MUX_Subtract23_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg311_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg22_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg338_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg338_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg279_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg118_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg285_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract23_0_impl_1_out);

   Delay1No197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_0_impl_1_out,
                 Y => Delay1No197_out);

Delay1No198_out_to_Subtract23_1_impl_parent_implementedSystem_port_0_cast <= Delay1No198_out;
Delay1No199_out_to_Subtract23_1_impl_parent_implementedSystem_port_1_cast <= Delay1No199_out;
   Subtract23_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract23_1_impl_out,
                 X => Delay1No198_out_to_Subtract23_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No199_out_to_Subtract23_1_impl_parent_implementedSystem_port_1_cast);

SharedReg321_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg321_out;
Delay4No23_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_2_cast <= Delay4No23_out;
SharedReg132_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg132_out;
SharedReg264_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg264_out;
SharedReg304_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg304_out;
SharedReg6_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg6_out;
SharedReg323_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg323_out;
   MUX_Subtract23_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg321_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No23_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg132_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg264_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg304_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg6_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg323_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract23_1_impl_0_out);

   Delay1No198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_1_impl_0_out,
                 Y => Delay1No198_out);

SharedReg337_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg337_out;
SharedReg289_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg289_out;
SharedReg123_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg123_out;
SharedReg288_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg288_out;
SharedReg315_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg315_out;
SharedReg22_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg22_out;
SharedReg339_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg339_out;
   MUX_Subtract23_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg337_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg289_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg123_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg288_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg315_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg22_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg339_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract23_1_impl_1_out);

   Delay1No199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_1_impl_1_out,
                 Y => Delay1No199_out);

Delay1No200_out_to_Product124_0_impl_parent_implementedSystem_port_0_cast <= Delay1No200_out;
Delay1No201_out_to_Product124_0_impl_parent_implementedSystem_port_1_cast <= Delay1No201_out;
   Product124_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product124_0_impl_out,
                 X => Delay1No200_out_to_Product124_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No201_out_to_Product124_0_impl_parent_implementedSystem_port_1_cast);

SharedReg406_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg406_out;
SharedReg436_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg436_out;
SharedReg400_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg400_out;
SharedReg427_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg427_out;
SharedReg425_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg425_out;
SharedReg402_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg402_out;
SharedReg392_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg392_out;
   MUX_Product124_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg406_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg436_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg400_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg427_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg425_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg402_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg392_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product124_0_impl_0_out);

   Delay1No200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_0_impl_0_out,
                 Y => Delay1No200_out);

SharedReg79_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg79_out;
SharedReg327_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg327_out;
SharedReg38_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg38_out;
SharedReg390_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg390_out;
SharedReg367_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg367_out;
SharedReg358_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg358_out;
SharedReg215_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg215_out;
   MUX_Product124_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg79_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg327_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg38_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg367_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg358_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg215_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product124_0_impl_1_out);

   Delay1No201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_0_impl_1_out,
                 Y => Delay1No201_out);

Delay1No202_out_to_Product124_1_impl_parent_implementedSystem_port_0_cast <= Delay1No202_out;
Delay1No203_out_to_Product124_1_impl_parent_implementedSystem_port_1_cast <= Delay1No203_out;
   Product124_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product124_1_impl_out,
                 X => Delay1No202_out_to_Product124_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No203_out_to_Product124_1_impl_parent_implementedSystem_port_1_cast);

SharedReg427_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg427_out;
SharedReg425_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg425_out;
SharedReg365_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg365_out;
SharedReg392_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg392_out;
SharedReg406_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg406_out;
SharedReg436_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg436_out;
SharedReg400_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg400_out;
   MUX_Product124_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg427_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg425_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg365_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg392_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg406_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg436_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg400_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product124_1_impl_0_out);

   Delay1No202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_1_impl_0_out,
                 Y => Delay1No202_out);

SharedReg388_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg388_out;
SharedReg355_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg355_out;
SharedReg417_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg417_out;
SharedReg218_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg218_out;
SharedReg82_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg82_out;
SharedReg332_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg332_out;
SharedReg41_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg41_out;
   MUX_Product124_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg388_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg355_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg417_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg218_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg82_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg332_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg41_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product124_1_impl_1_out);

   Delay1No203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_1_impl_1_out,
                 Y => Delay1No203_out);

Delay1No204_out_to_Product323_0_impl_parent_implementedSystem_port_0_cast <= Delay1No204_out;
Delay1No205_out_to_Product323_0_impl_parent_implementedSystem_port_1_cast <= Delay1No205_out;
   Product323_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product323_0_impl_out,
                 X => Delay1No204_out_to_Product323_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No205_out_to_Product323_0_impl_parent_implementedSystem_port_1_cast);

SharedReg393_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg393_out;
SharedReg327_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg327_out;
SharedReg400_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg400_out;
SharedReg431_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg431_out;
SharedReg429_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg429_out;
SharedReg402_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg402_out;
SharedReg392_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg392_out;
   MUX_Product323_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg393_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg327_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg400_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg431_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg429_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg402_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg392_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product323_0_impl_0_out);

   Delay1No204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_0_impl_0_out,
                 Y => Delay1No204_out);

SharedReg97_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg97_out;
SharedReg441_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg441_out;
SharedReg78_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg78_out;
SharedReg386_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg386_out;
SharedReg351_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg351_out;
SharedReg340_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg340_out;
SharedReg171_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg171_out;
   MUX_Product323_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg97_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg441_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg78_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg386_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg351_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg340_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg171_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product323_0_impl_1_out);

   Delay1No205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_0_impl_1_out,
                 Y => Delay1No205_out);

Delay1No206_out_to_Product323_1_impl_parent_implementedSystem_port_0_cast <= Delay1No206_out;
Delay1No207_out_to_Product323_1_impl_parent_implementedSystem_port_1_cast <= Delay1No207_out;
   Product323_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product323_1_impl_out,
                 X => Delay1No206_out_to_Product323_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No207_out_to_Product323_1_impl_parent_implementedSystem_port_1_cast);

SharedReg427_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg427_out;
SharedReg425_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg425_out;
SharedReg402_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg402_out;
SharedReg392_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg392_out;
SharedReg393_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg393_out;
SharedReg332_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg332_out;
SharedReg400_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg400_out;
   MUX_Product323_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg427_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg425_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg402_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg392_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg393_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg332_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg400_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product323_1_impl_0_out);

   Delay1No206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_1_impl_0_out,
                 Y => Delay1No206_out);

SharedReg391_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg370_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg370_out;
SharedReg362_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg362_out;
SharedReg175_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg175_out;
SharedReg101_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg101_out;
SharedReg441_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg441_out;
SharedReg81_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg81_out;
   MUX_Product323_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg370_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg362_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg175_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg101_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg441_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg81_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product323_1_impl_1_out);

   Delay1No207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_1_impl_1_out,
                 Y => Delay1No207_out);

Delay1No208_out_to_Product324_0_impl_parent_implementedSystem_port_0_cast <= Delay1No208_out;
Delay1No209_out_to_Product324_0_impl_parent_implementedSystem_port_1_cast <= Delay1No209_out;
   Product324_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product324_0_impl_out,
                 X => Delay1No208_out_to_Product324_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No209_out_to_Product324_0_impl_parent_implementedSystem_port_1_cast);

SharedReg97_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg97_out;
SharedReg86_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg86_out;
SharedReg413_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg413_out;
SharedReg390_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg390_out;
SharedReg367_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg367_out;
SharedReg415_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg415_out;
SharedReg405_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg405_out;
   MUX_Product324_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg97_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg86_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg413_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg367_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg415_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg405_out_to_MUX_Product324_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product324_0_impl_0_out);

   Delay1No208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product324_0_impl_0_out,
                 Y => Delay1No208_out);

SharedReg406_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg406_out;
SharedReg407_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg407_out;
SharedReg38_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg38_out;
SharedReg431_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg431_out;
SharedReg429_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg429_out;
SharedReg358_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg358_out;
SharedReg215_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg215_out;
   MUX_Product324_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg406_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg407_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg38_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg431_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg429_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg358_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg215_out_to_MUX_Product324_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product324_0_impl_1_out);

   Delay1No209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product324_0_impl_1_out,
                 Y => Delay1No209_out);

Delay1No210_out_to_Product324_1_impl_parent_implementedSystem_port_0_cast <= Delay1No210_out;
Delay1No211_out_to_Product324_1_impl_parent_implementedSystem_port_1_cast <= Delay1No211_out;
   Product324_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product324_1_impl_out,
                 X => Delay1No210_out_to_Product324_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No211_out_to_Product324_1_impl_parent_implementedSystem_port_1_cast);

SharedReg431_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg431_out;
SharedReg429_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg429_out;
SharedReg402_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg402_out;
SharedReg405_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg405_out;
SharedReg101_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg101_out;
SharedReg89_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg89_out;
SharedReg413_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg413_out;
   MUX_Product324_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg431_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg429_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg402_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg405_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg101_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg89_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg413_out_to_MUX_Product324_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product324_1_impl_0_out);

   Delay1No210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product324_1_impl_0_out,
                 Y => Delay1No210_out);

SharedReg388_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg388_out;
SharedReg355_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg355_out;
SharedReg345_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg345_out;
SharedReg218_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg218_out;
SharedReg406_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg406_out;
SharedReg407_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg407_out;
SharedReg41_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg41_out;
   MUX_Product324_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg388_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg355_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg345_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg218_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg406_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg407_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg41_out_to_MUX_Product324_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product324_1_impl_1_out);

   Delay1No211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product324_1_impl_1_out,
                 Y => Delay1No211_out);

Delay1No212_out_to_Product325_1_impl_parent_implementedSystem_port_0_cast <= Delay1No212_out;
Delay1No213_out_to_Product325_1_impl_parent_implementedSystem_port_1_cast <= Delay1No213_out;
   Product325_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product325_1_impl_out,
                 X => Delay1No212_out_to_Product325_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No213_out_to_Product325_1_impl_parent_implementedSystem_port_1_cast);

SharedReg391_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg370_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg370_out;
SharedReg415_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg415_out;
SharedReg175_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg175_out;
SharedReg393_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg393_out;
SharedReg436_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg436_out;
SharedReg81_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg81_out;
   MUX_Product325_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg370_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg415_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg175_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg393_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg436_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg81_out_to_MUX_Product325_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product325_1_impl_0_out);

   Delay1No212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product325_1_impl_0_out,
                 Y => Delay1No212_out);

SharedReg431_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg431_out;
SharedReg429_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg429_out;
SharedReg362_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg362_out;
SharedReg405_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg405_out;
SharedReg120_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg120_out;
SharedReg377_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg377_out;
SharedReg413_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg413_out;
   MUX_Product325_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg431_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg429_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg362_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg405_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg120_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg377_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg413_out_to_MUX_Product325_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product325_1_impl_1_out);

   Delay1No213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product325_1_impl_1_out,
                 Y => Delay1No213_out);

Delay1No214_out_to_Product55_0_impl_parent_implementedSystem_port_0_cast <= Delay1No214_out;
Delay1No215_out_to_Product55_0_impl_parent_implementedSystem_port_1_cast <= Delay1No215_out;
   Product55_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_0_impl_out,
                 X => Delay1No214_out_to_Product55_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No215_out_to_Product55_0_impl_parent_implementedSystem_port_1_cast);

SharedReg393_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg393_out;
SharedReg436_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg436_out;
SharedReg78_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg78_out;
SharedReg427_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg427_out;
SharedReg46_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg46_out;
SharedReg340_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg340_out;
SharedReg171_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg171_out;
   MUX_Product55_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg393_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg436_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg78_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg427_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg46_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg340_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg171_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product55_0_impl_0_out);

   Delay1No214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_0_impl_0_out,
                 Y => Delay1No214_out);

SharedReg115_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg115_out;
SharedReg373_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg373_out;
SharedReg413_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg413_out;
SharedReg372_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg372_out;
SharedReg416_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg416_out;
SharedReg415_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg415_out;
SharedReg405_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg405_out;
   MUX_Product55_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg115_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg373_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg413_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg372_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg416_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg415_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg405_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product55_0_impl_1_out);

   Delay1No215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_0_impl_1_out,
                 Y => Delay1No215_out);

Delay1No216_out_to_Product226_0_impl_parent_implementedSystem_port_0_cast <= Delay1No216_out;
Delay1No217_out_to_Product226_0_impl_parent_implementedSystem_port_1_cast <= Delay1No217_out;
   Product226_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product226_0_impl_out,
                 X => Delay1No216_out_to_Product226_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No217_out_to_Product226_0_impl_parent_implementedSystem_port_1_cast);

SharedReg115_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg115_out;
SharedReg441_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg441_out;
SharedReg426_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg426_out;
SharedReg427_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg427_out;
SharedReg403_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg403_out;
SharedReg402_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg402_out;
SharedReg448_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg448_out;
   MUX_Product226_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg115_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg441_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg426_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg427_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg403_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg402_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg448_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product226_0_impl_0_out);

   Delay1No216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_0_impl_0_out,
                 Y => Delay1No216_out);

SharedReg406_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg406_out;
SharedReg373_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg373_out;
SharedReg386_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg386_out;
SharedReg380_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg380_out;
SharedReg62_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg62_out;
SharedReg350_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg350_out;
SharedReg187_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg187_out;
   MUX_Product226_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg406_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg373_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg386_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg380_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg62_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg350_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg187_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product226_0_impl_1_out);

   Delay1No217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_0_impl_1_out,
                 Y => Delay1No217_out);

Delay1No218_out_to_Product226_1_impl_parent_implementedSystem_port_0_cast <= Delay1No218_out;
Delay1No219_out_to_Product226_1_impl_parent_implementedSystem_port_1_cast <= Delay1No219_out;
   Product226_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product226_1_impl_out,
                 X => Delay1No218_out_to_Product226_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No219_out_to_Product226_1_impl_parent_implementedSystem_port_1_cast);

SharedReg427_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg427_out;
SharedReg51_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg51_out;
SharedReg345_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg345_out;
SharedReg448_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg448_out;
SharedReg120_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg120_out;
SharedReg441_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg441_out;
SharedReg426_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg426_out;
   MUX_Product226_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg427_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg51_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg345_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg448_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg120_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg441_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg426_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product226_1_impl_0_out);

   Delay1No218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_1_impl_0_out,
                 Y => Delay1No218_out);

SharedReg376_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg376_out;
SharedReg416_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg416_out;
SharedReg415_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg415_out;
SharedReg191_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg191_out;
SharedReg406_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg406_out;
SharedReg377_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg377_out;
SharedReg388_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg388_out;
   MUX_Product226_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg376_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg416_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg415_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg191_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg406_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg377_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg388_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product226_1_impl_1_out);

   Delay1No219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_1_impl_1_out,
                 Y => Delay1No219_out);

Delay1No220_out_to_Product130_1_impl_parent_implementedSystem_port_0_cast <= Delay1No220_out;
Delay1No221_out_to_Product130_1_impl_parent_implementedSystem_port_1_cast <= Delay1No221_out;
   Product130_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product130_1_impl_out,
                 X => Delay1No220_out_to_Product130_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No221_out_to_Product130_1_impl_parent_implementedSystem_port_1_cast);

SharedReg427_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg427_out;
SharedReg403_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg403_out;
SharedReg402_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg402_out;
SharedReg448_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg448_out;
SharedReg393_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg393_out;
SharedReg394_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg394_out;
SharedReg426_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg426_out;
   MUX_Product130_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg427_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg403_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg402_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg448_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg393_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg394_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg426_out_to_MUX_Product130_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product130_1_impl_0_out);

   Delay1No220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product130_1_impl_0_out,
                 Y => Delay1No220_out);

SharedReg383_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg383_out;
SharedReg65_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg65_out;
SharedReg354_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg354_out;
SharedReg236_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg236_out;
SharedReg142_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg142_out;
SharedReg94_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg94_out;
SharedReg391_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg391_out;
   MUX_Product130_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg383_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg65_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg354_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg236_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg142_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg94_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg391_out_to_MUX_Product130_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product130_1_impl_1_out);

   Delay1No221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product130_1_impl_1_out,
                 Y => Delay1No221_out);

Delay1No222_out_to_Product329_0_impl_parent_implementedSystem_port_0_cast <= Delay1No222_out;
Delay1No223_out_to_Product329_0_impl_parent_implementedSystem_port_1_cast <= Delay1No223_out;
   Product329_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product329_0_impl_out,
                 X => Delay1No222_out_to_Product329_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No223_out_to_Product329_0_impl_parent_implementedSystem_port_1_cast);

SharedReg393_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg393_out;
SharedReg394_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg394_out;
SharedReg426_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg426_out;
SharedReg431_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg431_out;
SharedReg62_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg62_out;
SharedReg402_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg402_out;
SharedReg448_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg448_out;
   MUX_Product329_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg393_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg394_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg426_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg431_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg62_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg402_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg448_out_to_MUX_Product329_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product329_0_impl_0_out);

   Delay1No222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product329_0_impl_0_out,
                 Y => Delay1No222_out);

SharedReg137_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg137_out;
SharedReg91_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg91_out;
SharedReg390_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg372_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg372_out;
SharedReg416_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg416_out;
SharedReg366_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg366_out;
SharedReg233_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg233_out;
   MUX_Product329_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg137_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg91_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg372_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg416_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg366_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg233_out_to_MUX_Product329_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product329_0_impl_1_out);

   Delay1No223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product329_0_impl_1_out,
                 Y => Delay1No223_out);

Delay1No224_out_to_Product329_1_impl_parent_implementedSystem_port_0_cast <= Delay1No224_out;
Delay1No225_out_to_Product329_1_impl_parent_implementedSystem_port_1_cast <= Delay1No225_out;
   Product329_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product329_1_impl_out,
                 X => Delay1No224_out_to_Product329_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No225_out_to_Product329_1_impl_parent_implementedSystem_port_1_cast);

SharedReg431_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg431_out;
SharedReg65_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg65_out;
SharedReg402_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg402_out;
SharedReg449_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg449_out;
SharedReg393_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg393_out;
SharedReg407_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg407_out;
SharedReg430_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg430_out;
   MUX_Product329_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg431_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg65_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg402_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg449_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg393_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg407_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg430_out_to_MUX_Product329_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product329_1_impl_0_out);

   Delay1No224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product329_1_impl_0_out,
                 Y => Delay1No224_out);

SharedReg376_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg376_out;
SharedReg416_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg416_out;
SharedReg369_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg369_out;
SharedReg191_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg191_out;
SharedReg152_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg152_out;
SharedReg94_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg94_out;
SharedReg388_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg388_out;
   MUX_Product329_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg376_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg416_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg369_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg191_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg152_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg94_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg388_out_to_MUX_Product329_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product329_1_impl_1_out);

   Delay1No225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product329_1_impl_1_out,
                 Y => Delay1No225_out);

Delay1No226_out_to_Subtract30_0_impl_parent_implementedSystem_port_0_cast <= Delay1No226_out;
Delay1No227_out_to_Subtract30_0_impl_parent_implementedSystem_port_1_cast <= Delay1No227_out;
   Subtract30_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract30_0_impl_out,
                 X => Delay1No226_out_to_Subtract30_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No227_out_to_Subtract30_0_impl_parent_implementedSystem_port_1_cast);

SharedReg317_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg317_out;
SharedReg7_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg7_out;
SharedReg136_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg136_out;
SharedReg254_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg254_out;
SharedReg206_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg206_out;
SharedReg97_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg97_out;
SharedReg116_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg116_out;
   MUX_Subtract30_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg317_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg136_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg254_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg206_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg97_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg116_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract30_0_impl_0_out);

   Delay1No226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_0_impl_0_out,
                 Y => Delay1No226_out);

SharedReg336_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg336_out;
SharedReg23_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg23_out;
SharedReg146_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg146_out;
SharedReg341_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg341_out;
Delay4No32_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_5_cast <= Delay4No32_out;
SharedReg129_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg129_out;
SharedReg140_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg140_out;
   MUX_Subtract30_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg336_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg23_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg146_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg341_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay4No32_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg129_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg140_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract30_0_impl_1_out);

   Delay1No227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_0_impl_1_out,
                 Y => Delay1No227_out);

Delay1No228_out_to_Subtract30_1_impl_parent_implementedSystem_port_0_cast <= Delay1No228_out;
Delay1No229_out_to_Subtract30_1_impl_parent_implementedSystem_port_1_cast <= Delay1No229_out;
   Subtract30_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract30_1_impl_out,
                 X => Delay1No228_out_to_Subtract30_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No229_out_to_Subtract30_1_impl_parent_implementedSystem_port_1_cast);

SharedReg258_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg258_out;
SharedReg214_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg214_out;
SharedReg101_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg101_out;
SharedReg121_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg121_out;
SharedReg321_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg321_out;
SharedReg7_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg7_out;
SharedReg141_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg141_out;
   MUX_Subtract30_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg258_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg214_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg101_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg121_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg321_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg7_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg141_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract30_1_impl_0_out);

   Delay1No228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_1_impl_0_out,
                 Y => Delay1No228_out);

SharedReg346_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg346_out;
Delay4No33_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_2_cast <= Delay4No33_out;
SharedReg135_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg135_out;
SharedReg145_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg145_out;
SharedReg337_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg337_out;
SharedReg23_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg23_out;
SharedReg151_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg151_out;
   MUX_Subtract30_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg346_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No33_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg135_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg145_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg337_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg23_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg151_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract30_1_impl_1_out);

   Delay1No229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_1_impl_1_out,
                 Y => Delay1No229_out);

Delay1No230_out_to_Product132_0_impl_parent_implementedSystem_port_0_cast <= Delay1No230_out;
Delay1No231_out_to_Product132_0_impl_parent_implementedSystem_port_1_cast <= Delay1No231_out;
   Product132_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product132_0_impl_out,
                 X => Delay1No230_out_to_Product132_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No231_out_to_Product132_0_impl_parent_implementedSystem_port_1_cast);

SharedReg393_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg393_out;
SharedReg407_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg407_out;
SharedReg430_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg430_out;
SharedReg380_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg380_out;
SharedReg403_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg403_out;
SharedReg415_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg415_out;
SharedReg449_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg449_out;
   MUX_Product132_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg393_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg407_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg430_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg380_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg403_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg415_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg449_out_to_MUX_Product132_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product132_0_impl_0_out);

   Delay1No230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product132_0_impl_0_out,
                 Y => Delay1No230_out);

SharedReg147_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg147_out;
SharedReg91_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg91_out;
SharedReg386_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg386_out;
SharedReg431_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg431_out;
SharedReg343_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg343_out;
SharedReg350_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg350_out;
SharedReg187_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg187_out;
   MUX_Product132_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg147_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg91_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg386_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg431_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg343_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg350_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg187_out_to_MUX_Product132_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product132_0_impl_1_out);

   Delay1No231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product132_0_impl_1_out,
                 Y => Delay1No231_out);

Delay1No232_out_to_Product132_1_impl_parent_implementedSystem_port_0_cast <= Delay1No232_out;
Delay1No233_out_to_Product132_1_impl_parent_implementedSystem_port_1_cast <= Delay1No233_out;
   Product132_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product132_1_impl_out,
                 X => Delay1No232_out_to_Product132_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No233_out_to_Product132_1_impl_parent_implementedSystem_port_1_cast);

SharedReg383_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg383_out;
SharedReg403_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg403_out;
SharedReg415_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg415_out;
SharedReg236_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg236_out;
SharedReg406_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg406_out;
SharedReg394_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg394_out;
SharedReg391_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg391_out;
   MUX_Product132_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg383_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg403_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg415_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg236_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg406_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg394_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg391_out_to_MUX_Product132_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product132_1_impl_0_out);

   Delay1No232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product132_1_impl_0_out,
                 Y => Delay1No232_out);

SharedReg431_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg431_out;
SharedReg348_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg348_out;
SharedReg354_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg354_out;
SharedReg449_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg449_out;
SharedReg142_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg142_out;
SharedReg111_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg111_out;
SharedReg430_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg430_out;
   MUX_Product132_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg431_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg348_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg354_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg449_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg142_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg111_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg430_out_to_MUX_Product132_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product132_1_impl_1_out);

   Delay1No233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product132_1_impl_1_out,
                 Y => Delay1No233_out);

Delay1No234_out_to_Product331_0_impl_parent_implementedSystem_port_0_cast <= Delay1No234_out;
Delay1No235_out_to_Product331_0_impl_parent_implementedSystem_port_1_cast <= Delay1No235_out;
   Product331_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product331_0_impl_out,
                 X => Delay1No234_out_to_Product331_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No235_out_to_Product331_0_impl_parent_implementedSystem_port_1_cast);

SharedReg406_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg406_out;
SharedReg394_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg394_out;
SharedReg390_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg408_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg408_out;
SharedReg343_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg343_out;
SharedReg366_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg366_out;
SharedReg233_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg233_out;
   MUX_Product331_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg406_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg394_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg408_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg343_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg366_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg233_out_to_MUX_Product331_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product331_0_impl_0_out);

   Delay1No234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product331_0_impl_0_out,
                 Y => Delay1No234_out);

SharedReg137_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg137_out;
SharedReg106_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg106_out;
SharedReg430_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg430_out;
Delay5No8_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_4_cast <= Delay5No8_out;
SharedReg416_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg416_out;
SharedReg415_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg415_out;
SharedReg449_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg449_out;
   MUX_Product331_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg137_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg106_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg430_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay5No8_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg416_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg415_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg449_out_to_MUX_Product331_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Product331_0_impl_1_out);

   Delay1No235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product331_0_impl_1_out,
                 Y => Delay1No235_out);

Delay1No236_out_to_Product331_1_impl_parent_implementedSystem_port_0_cast <= Delay1No236_out;
Delay1No237_out_to_Product331_1_impl_parent_implementedSystem_port_1_cast <= Delay1No237_out;
   Product331_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product331_1_impl_out,
                 X => Delay1No236_out_to_Product331_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No237_out_to_Product331_1_impl_parent_implementedSystem_port_1_cast);

SharedReg152_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg152_out;
SharedReg348_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg348_out;
SharedReg369_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg369_out;
SharedReg407_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg407_out;
SharedReg395_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg395_out;
SharedReg408_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg408_out;
   MUX_Product331_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg152_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg348_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg369_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg407_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg395_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg408_out_to_MUX_Product331_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => MUX_Product331_1_impl_0_LUT_out,
                 oMux => MUX_Product331_1_impl_0_out);

   Delay1No236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product331_1_impl_0_out,
                 Y => Delay1No236_out);

SharedReg111_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg77_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg77_out;
Delay5No9_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_3_cast <= Delay5No9_out;
SharedReg416_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg416_out;
SharedReg415_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg415_out;
SharedReg406_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg406_out;
   MUX_Product331_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg77_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay5No9_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg416_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg415_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg406_out_to_MUX_Product331_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => MUX_Product331_1_impl_1_LUT_out,
                 oMux => MUX_Product331_1_impl_1_out);

   Delay1No237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product331_1_impl_1_out,
                 Y => Delay1No237_out);

Delay1No238_out_to_Subtract42_0_impl_parent_implementedSystem_port_0_cast <= Delay1No238_out;
Delay1No239_out_to_Subtract42_0_impl_parent_implementedSystem_port_1_cast <= Delay1No239_out;
   Subtract42_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract42_0_impl_out,
                 X => Delay1No238_out_to_Subtract42_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No239_out_to_Subtract42_0_impl_parent_implementedSystem_port_1_cast);

SharedReg96_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg96_out;
SharedReg9_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg9_out;
SharedReg137_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg137_out;
SharedReg116_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg116_out;
SharedReg324_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg324_out;
SharedReg99_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg99_out;
SharedReg302_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg302_out;
   MUX_Subtract42_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg96_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg9_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg137_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg116_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg324_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg99_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg302_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract42_0_impl_0_out);

   Delay1No238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_0_impl_0_out,
                 Y => Delay1No238_out);

SharedReg104_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg104_out;
SharedReg25_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg25_out;
SharedReg96_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg96_out;
SharedReg125_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg125_out;
SharedReg165_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg165_out;
SharedReg146_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg146_out;
SharedReg317_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg317_out;
   MUX_Subtract42_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg104_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg25_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg96_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg125_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg165_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg146_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg317_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract42_0_impl_1_out);

   Delay1No239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_0_impl_1_out,
                 Y => Delay1No239_out);

Delay1No240_out_to_Subtract42_1_impl_parent_implementedSystem_port_0_cast <= Delay1No240_out;
Delay1No241_out_to_Subtract42_1_impl_parent_implementedSystem_port_1_cast <= Delay1No241_out;
   Subtract42_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract42_1_impl_out,
                 X => Delay1No240_out_to_Subtract42_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No241_out_to_Subtract42_1_impl_parent_implementedSystem_port_1_cast);

SharedReg121_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg121_out;
SharedReg323_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg323_out;
SharedReg103_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg103_out;
SharedReg304_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg304_out;
SharedReg100_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg100_out;
SharedReg9_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg9_out;
SharedReg142_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg142_out;
   MUX_Subtract42_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg121_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg323_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg103_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg304_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg100_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg9_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg142_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract42_1_impl_0_out);

   Delay1No240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_1_impl_0_out,
                 Y => Delay1No240_out);

SharedReg131_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg339_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg339_out;
SharedReg151_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg151_out;
SharedReg315_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg315_out;
SharedReg109_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg109_out;
SharedReg25_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg100_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg100_out;
   MUX_Subtract42_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg339_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg151_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg315_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg109_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg25_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg100_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract42_1_impl_1_out);

   Delay1No241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_1_impl_1_out,
                 Y => Delay1No241_out);

Delay1No242_out_to_Subtract44_0_impl_parent_implementedSystem_port_0_cast <= Delay1No242_out;
Delay1No243_out_to_Subtract44_0_impl_parent_implementedSystem_port_1_cast <= Delay1No243_out;
   Subtract44_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract44_0_impl_out,
                 X => Delay1No242_out_to_Subtract44_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No243_out_to_Subtract44_0_impl_parent_implementedSystem_port_1_cast);

SharedReg187_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg187_out;
SharedReg10_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg10_out;
SharedReg291_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg291_out;
SharedReg255_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg255_out;
SharedReg173_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg173_out;
SharedReg217_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg217_out;
SharedReg319_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg319_out;
   MUX_Subtract44_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg187_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg291_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg255_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg173_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg217_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg319_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract44_0_impl_0_out);

   Delay1No242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_0_impl_0_out,
                 Y => Delay1No242_out);

SharedReg233_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg233_out;
SharedReg26_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg26_out;
SharedReg254_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg254_out;
SharedReg344_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg344_out;
SharedReg366_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg366_out;
SharedReg215_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg215_out;
SharedReg338_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg338_out;
   MUX_Subtract44_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg233_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg26_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg254_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg344_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg366_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg215_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg338_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract44_0_impl_1_out);

   Delay1No243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_0_impl_1_out,
                 Y => Delay1No243_out);

Delay1No244_out_to_Subtract44_1_impl_parent_implementedSystem_port_0_cast <= Delay1No244_out;
Delay1No245_out_to_Subtract44_1_impl_parent_implementedSystem_port_1_cast <= Delay1No245_out;
   Subtract44_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract44_1_impl_out,
                 X => Delay1No244_out_to_Subtract44_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No245_out_to_Subtract44_1_impl_parent_implementedSystem_port_1_cast);

SharedReg259_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg259_out;
SharedReg177_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg177_out;
SharedReg220_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg220_out;
SharedReg321_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg321_out;
SharedReg191_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg191_out;
SharedReg10_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg10_out;
SharedReg297_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg297_out;
   MUX_Subtract44_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg259_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg177_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg220_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg321_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg191_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg10_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg297_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract44_1_impl_0_out);

   Delay1No244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_1_impl_0_out,
                 Y => Delay1No244_out);

SharedReg349_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg349_out;
SharedReg369_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg369_out;
SharedReg218_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg218_out;
SharedReg337_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg337_out;
SharedReg236_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg236_out;
SharedReg26_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg26_out;
SharedReg258_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg258_out;
   MUX_Subtract44_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg349_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg369_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg218_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg337_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg236_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg26_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg258_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract44_1_impl_1_out);

   Delay1No245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_1_impl_1_out,
                 Y => Delay1No245_out);

Delay1No246_out_to_Subtract45_0_impl_parent_implementedSystem_port_0_cast <= Delay1No246_out;
Delay1No247_out_to_Subtract45_0_impl_parent_implementedSystem_port_1_cast <= Delay1No247_out;
   Subtract45_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract45_0_impl_out,
                 X => Delay1No246_out_to_Subtract45_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No247_out_to_Subtract45_0_impl_parent_implementedSystem_port_1_cast);

SharedReg215_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg215_out;
SharedReg8_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
SharedReg270_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg270_out;
SharedReg80_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg80_out;
SharedReg328_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg328_out;
SharedReg338_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg338_out;
SharedReg234_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg234_out;
   MUX_Subtract45_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg215_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg270_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg80_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg328_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg338_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg234_out_to_MUX_Subtract45_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract45_0_impl_0_out);

   Delay1No246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract45_0_impl_0_out,
                 Y => Delay1No246_out);

SharedReg171_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg171_out;
SharedReg24_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg233_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg233_out;
SharedReg106_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg106_out;
SharedReg272_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg272_out;
SharedReg320_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg320_out;
SharedReg295_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg295_out;
   MUX_Subtract45_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg171_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg233_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg106_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg272_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg320_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg295_out_to_MUX_Subtract45_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract45_0_impl_1_out);

   Delay1No247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract45_0_impl_1_out,
                 Y => Delay1No247_out);

Delay1No248_out_to_Subtract45_1_impl_parent_implementedSystem_port_0_cast <= Delay1No248_out;
Delay1No249_out_to_Subtract45_1_impl_parent_implementedSystem_port_1_cast <= Delay1No249_out;
   Subtract45_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract45_1_impl_out,
                 X => Delay1No248_out_to_Subtract45_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No249_out_to_Subtract45_1_impl_parent_implementedSystem_port_1_cast);

SharedReg83_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg83_out;
SharedReg333_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg333_out;
SharedReg337_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg337_out;
SharedReg237_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg237_out;
SharedReg218_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg218_out;
SharedReg8_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg8_out;
SharedReg274_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg274_out;
   MUX_Subtract45_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg83_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg333_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg337_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg237_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg218_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg8_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg274_out_to_MUX_Subtract45_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract45_1_impl_0_out);

   Delay1No248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract45_1_impl_0_out,
                 Y => Delay1No248_out);

SharedReg111_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg276_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg276_out;
SharedReg322_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg322_out;
SharedReg301_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg301_out;
SharedReg175_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg175_out;
SharedReg24_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg24_out;
SharedReg236_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg236_out;
   MUX_Subtract45_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg276_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg322_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg301_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg24_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg236_out_to_MUX_Subtract45_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract45_1_impl_1_out);

   Delay1No249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract45_1_impl_1_out,
                 Y => Delay1No249_out);

Delay1No250_out_to_Subtract46_0_impl_parent_implementedSystem_port_0_cast <= Delay1No250_out;
Delay1No251_out_to_Subtract46_0_impl_parent_implementedSystem_port_1_cast <= Delay1No251_out;
   Subtract46_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract46_0_impl_out,
                 X => Delay1No250_out_to_Subtract46_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No251_out_to_Subtract46_0_impl_parent_implementedSystem_port_1_cast);

SharedReg86_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg86_out;
SharedReg11_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg11_out;
SharedReg147_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg147_out;
SharedReg126_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg126_out;
SharedReg235_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg235_out;
SharedReg92_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg92_out;
SharedReg165_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg165_out;
   MUX_Subtract46_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg86_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg11_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg147_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg126_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg235_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg92_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg165_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract46_0_impl_0_out);

   Delay1No250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_0_impl_0_out,
                 Y => Delay1No250_out);

SharedReg114_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg114_out;
SharedReg27_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg27_out;
SharedReg104_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg104_out;
SharedReg139_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg139_out;
SharedReg292_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg292_out;
SharedReg72_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg72_out;
SharedReg287_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg287_out;
   MUX_Subtract46_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg114_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg104_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg139_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg292_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg72_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg287_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract46_0_impl_1_out);

   Delay1No251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_0_impl_1_out,
                 Y => Delay1No251_out);

Delay1No252_out_to_Subtract46_1_impl_parent_implementedSystem_port_0_cast <= Delay1No252_out;
Delay1No253_out_to_Subtract46_1_impl_parent_implementedSystem_port_1_cast <= Delay1No253_out;
   Subtract46_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract46_1_impl_out,
                 X => Delay1No252_out_to_Subtract46_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No253_out_to_Subtract46_1_impl_parent_implementedSystem_port_1_cast);

SharedReg132_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg132_out;
SharedReg238_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg238_out;
SharedReg95_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg95_out;
SharedReg339_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg339_out;
SharedReg89_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg89_out;
SharedReg11_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg11_out;
SharedReg152_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg152_out;
   MUX_Subtract46_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg132_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg238_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg95_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg339_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg89_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg11_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg152_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract46_1_impl_0_out);

   Delay1No252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_1_impl_0_out,
                 Y => Delay1No252_out);

SharedReg144_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg144_out;
SharedReg298_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg298_out;
SharedReg75_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg75_out;
SharedReg289_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg289_out;
SharedReg119_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg119_out;
SharedReg27_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg27_out;
SharedReg109_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg109_out;
   MUX_Subtract46_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg144_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg298_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg75_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg289_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg119_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg27_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg109_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract46_1_impl_1_out);

   Delay1No253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_1_impl_1_out,
                 Y => Delay1No253_out);

Delay1No254_out_to_Subtract57_0_impl_parent_implementedSystem_port_0_cast <= Delay1No254_out;
Delay1No255_out_to_Subtract57_0_impl_parent_implementedSystem_port_1_cast <= Delay1No255_out;
   Subtract57_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract57_0_impl_out,
                 X => Delay1No254_out_to_Subtract57_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No255_out_to_Subtract57_0_impl_parent_implementedSystem_port_1_cast);

SharedReg254_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg254_out;
SharedReg12_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg12_out;
SharedReg215_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg215_out;
SharedReg172_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg172_out;
SharedReg172_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg172_out;
SharedReg216_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg216_out;
SharedReg174_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg174_out;
   MUX_Subtract57_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg254_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg215_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg172_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg172_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg216_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg174_out_to_MUX_Subtract57_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract57_0_impl_0_out);

   Delay1No254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract57_0_impl_0_out,
                 Y => Delay1No254_out);

SharedReg256_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg256_out;
SharedReg28_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg28_out;
SharedReg269_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg269_out;
SharedReg269_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg269_out;
SharedReg215_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg215_out;
SharedReg187_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg187_out;
SharedReg190_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg190_out;
   MUX_Subtract57_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg256_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg28_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg269_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg269_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg215_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg187_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg190_out_to_MUX_Subtract57_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract57_0_impl_1_out);

   Delay1No255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract57_0_impl_1_out,
                 Y => Delay1No255_out);

Delay1No256_out_to_Subtract57_1_impl_parent_implementedSystem_port_0_cast <= Delay1No256_out;
Delay1No257_out_to_Subtract57_1_impl_parent_implementedSystem_port_1_cast <= Delay1No257_out;
   Subtract57_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract57_1_impl_out,
                 X => Delay1No256_out_to_Subtract57_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No257_out_to_Subtract57_1_impl_parent_implementedSystem_port_1_cast);

SharedReg176_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg176_out;
SharedReg176_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg176_out;
SharedReg219_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg219_out;
SharedReg178_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg178_out;
SharedReg258_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg258_out;
SharedReg12_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg12_out;
SharedReg218_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg218_out;
   MUX_Subtract57_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg176_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg176_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg219_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg178_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg258_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg12_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg218_out_to_MUX_Subtract57_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract57_1_impl_0_out);

   Delay1No256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract57_1_impl_0_out,
                 Y => Delay1No256_out);

SharedReg273_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg273_out;
SharedReg218_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg218_out;
SharedReg191_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg191_out;
SharedReg194_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg194_out;
SharedReg260_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg260_out;
SharedReg28_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg28_out;
SharedReg273_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg273_out;
   MUX_Subtract57_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg273_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg218_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg191_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg194_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg260_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg28_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg273_out_to_MUX_Subtract57_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract57_1_impl_1_out);

   Delay1No257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract57_1_impl_1_out,
                 Y => Delay1No257_out);

Delay1No258_out_to_Subtract117_0_impl_parent_implementedSystem_port_0_cast <= Delay1No258_out;
Delay1No259_out_to_Subtract117_0_impl_parent_implementedSystem_port_1_cast <= Delay1No259_out;
   Subtract117_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract117_0_impl_out,
                 X => Delay1No258_out_to_Subtract117_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No259_out_to_Subtract117_0_impl_parent_implementedSystem_port_1_cast);

SharedReg124_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg124_out;
SharedReg13_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg90_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg90_out;
SharedReg85_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg85_out;
SharedReg97_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg97_out;
SharedReg91_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg91_out;
SharedReg189_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg189_out;
   MUX_Subtract117_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg124_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg90_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg85_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg97_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg91_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg189_out_to_MUX_Subtract117_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract117_0_impl_0_out);

   Delay1No258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract117_0_impl_0_out,
                 Y => Delay1No258_out);

SharedReg107_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg107_out;
SharedReg29_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg29_out;
SharedReg114_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg114_out;
SharedReg136_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg136_out;
SharedReg78_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg78_out;
SharedReg90_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg90_out;
SharedReg257_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg257_out;
   MUX_Subtract117_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg107_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg114_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg136_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg78_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg90_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg257_out_to_MUX_Subtract117_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract117_0_impl_1_out);

   Delay1No259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract117_0_impl_1_out,
                 Y => Delay1No259_out);

Delay1No260_out_to_Subtract117_1_impl_parent_implementedSystem_port_0_cast <= Delay1No260_out;
Delay1No261_out_to_Subtract117_1_impl_parent_implementedSystem_port_1_cast <= Delay1No261_out;
   Subtract117_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract117_1_impl_out,
                 X => Delay1No260_out_to_Subtract117_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No261_out_to_Subtract117_1_impl_parent_implementedSystem_port_1_cast);

SharedReg88_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg88_out;
SharedReg101_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg101_out;
SharedReg94_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg94_out;
SharedReg193_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg193_out;
SharedReg130_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg130_out;
SharedReg13_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg13_out;
SharedReg93_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg93_out;
   MUX_Subtract117_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg88_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg101_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg94_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg193_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg130_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg13_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg93_out_to_MUX_Subtract117_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract117_1_impl_0_out);

   Delay1No260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract117_1_impl_0_out,
                 Y => Delay1No260_out);

SharedReg141_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg141_out;
SharedReg81_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg81_out;
SharedReg93_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg93_out;
SharedReg261_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg261_out;
SharedReg112_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg112_out;
SharedReg29_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg29_out;
SharedReg119_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg119_out;
   MUX_Subtract117_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg141_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg81_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg93_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg261_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg112_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg29_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg119_out_to_MUX_Subtract117_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract117_1_impl_1_out);

   Delay1No261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract117_1_impl_1_out,
                 Y => Delay1No261_out);

Delay1No262_out_to_Subtract61_0_impl_parent_implementedSystem_port_0_cast <= Delay1No262_out;
Delay1No263_out_to_Subtract61_0_impl_parent_implementedSystem_port_1_cast <= Delay1No263_out;
   Subtract61_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract61_0_impl_out,
                 X => Delay1No262_out_to_Subtract61_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No263_out_to_Subtract61_0_impl_parent_implementedSystem_port_1_cast);

SharedReg269_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg269_out;
SharedReg14_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg14_out;
SharedReg292_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg292_out;
SharedReg188_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg188_out;
SharedReg188_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg188_out;
SharedReg234_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg234_out;
SharedReg91_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg91_out;
   MUX_Subtract61_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg269_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg14_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg292_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg188_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg188_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg234_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg91_out_to_MUX_Subtract61_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract61_0_impl_0_out);

   Delay1No262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract61_0_impl_0_out,
                 Y => Delay1No262_out);

SharedReg293_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg293_out;
SharedReg30_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg30_out;
SharedReg353_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg353_out;
SharedReg358_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg358_out;
SharedReg171_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg171_out;
SharedReg233_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg233_out;
SharedReg108_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg108_out;
   MUX_Subtract61_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg293_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg353_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg358_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg171_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg233_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg108_out_to_MUX_Subtract61_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract61_0_impl_1_out);

   Delay1No263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract61_0_impl_1_out,
                 Y => Delay1No263_out);

Delay1No264_out_to_Subtract61_1_impl_parent_implementedSystem_port_0_cast <= Delay1No264_out;
Delay1No265_out_to_Subtract61_1_impl_parent_implementedSystem_port_1_cast <= Delay1No265_out;
   Subtract61_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract61_1_impl_out,
                 X => Delay1No264_out_to_Subtract61_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No265_out_to_Subtract61_1_impl_parent_implementedSystem_port_1_cast);

SharedReg192_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg192_out;
SharedReg192_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg192_out;
SharedReg237_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg237_out;
SharedReg94_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg94_out;
SharedReg273_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg273_out;
SharedReg14_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg14_out;
SharedReg298_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg298_out;
   MUX_Subtract61_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg192_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg192_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg237_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg94_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg273_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg14_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg298_out_to_MUX_Subtract61_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract61_1_impl_0_out);

   Delay1No264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract61_1_impl_0_out,
                 Y => Delay1No264_out);

SharedReg362_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg362_out;
SharedReg175_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg175_out;
SharedReg236_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg236_out;
SharedReg113_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg113_out;
SharedReg299_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg299_out;
SharedReg30_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg30_out;
SharedReg357_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg357_out;
   MUX_Subtract61_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg362_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg175_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg236_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg113_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg299_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg30_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg357_out_to_MUX_Subtract61_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract61_1_impl_1_out);

   Delay1No265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract61_1_impl_1_out,
                 Y => Delay1No265_out);

Delay1No266_out_to_Subtract121_0_impl_parent_implementedSystem_port_0_cast <= Delay1No266_out;
Delay1No267_out_to_Subtract121_0_impl_parent_implementedSystem_port_1_cast <= Delay1No267_out;
   Subtract121_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract121_0_impl_out,
                 X => Delay1No266_out_to_Subtract121_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No267_out_to_Subtract121_0_impl_parent_implementedSystem_port_1_cast);

SharedReg136_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg15_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg148_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg148_out;
SharedReg86_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg86_out;
SharedReg105_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg105_out;
SharedReg116_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg116_out;
SharedReg271_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg271_out;
   MUX_Subtract121_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg148_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg86_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg105_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg116_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg271_out_to_MUX_Subtract121_0_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract121_0_impl_0_out);

   Delay1No266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract121_0_impl_0_out,
                 Y => Delay1No266_out);

SharedReg127_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg127_out;
SharedReg31_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg31_out;
SharedReg150_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg150_out;
SharedReg146_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg146_out;
SharedReg84_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg84_out;
SharedReg96_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg96_out;
SharedReg330_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg330_out;
   MUX_Subtract121_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg150_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg146_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg84_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg96_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg330_out_to_MUX_Subtract121_0_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract121_0_impl_1_out);

   Delay1No267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract121_0_impl_1_out,
                 Y => Delay1No267_out);

Delay1No268_out_to_Subtract121_1_impl_parent_implementedSystem_port_0_cast <= Delay1No268_out;
Delay1No269_out_to_Subtract121_1_impl_parent_implementedSystem_port_1_cast <= Delay1No269_out;
   Subtract121_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract121_1_impl_out,
                 X => Delay1No268_out_to_Subtract121_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No269_out_to_Subtract121_1_impl_parent_implementedSystem_port_1_cast);

SharedReg89_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg89_out;
SharedReg110_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg110_out;
SharedReg121_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg121_out;
SharedReg275_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg275_out;
SharedReg141_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg141_out;
SharedReg15_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg15_out;
SharedReg153_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg153_out;
   MUX_Subtract121_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg89_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg110_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg121_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg275_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg141_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg15_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg153_out_to_MUX_Subtract121_1_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract121_1_impl_0_out);

   Delay1No268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract121_1_impl_0_out,
                 Y => Delay1No268_out);

SharedReg151_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg151_out;
SharedReg87_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg87_out;
SharedReg100_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg100_out;
SharedReg335_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg335_out;
SharedReg133_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg133_out;
SharedReg31_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg31_out;
SharedReg155_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg155_out;
   MUX_Subtract121_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg151_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg87_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg100_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg335_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg133_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg31_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg155_out_to_MUX_Subtract121_1_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => ModCount71_out,
                 oMux => MUX_Subtract121_1_impl_1_out);

   Delay1No269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract121_1_impl_1_out,
                 Y => Delay1No269_out);
   Constant2_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant2_0_impl_out);
   Constant11_0_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant11_0_impl_out);
   Constant4_0_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant4_0_impl_out);
   Constant13_0_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant13_0_impl_out);
   Constant5_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant5_0_impl_out);
   Constant14_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant14_0_impl_out);
   Constant6_0_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant6_0_impl_out);
   Constant15_0_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant15_0_impl_out);
   Constant7_0_impl_instance: Constant_float_8_23_cosn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant7_0_impl_out);
   Constant16_0_impl_instance: Constant_float_8_23_sinn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant16_0_impl_out);
   Constant8_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant8_0_impl_out);
   Constant17_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant17_0_impl_out);
   Constant9_0_impl_instance: Constant_float_8_23_cosn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant9_0_impl_out);
   Constant18_0_impl_instance: Constant_float_8_23_sinn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant18_0_impl_out);
   Constant_0_impl_instance: Constant_float_8_23_cosnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);
   Constant1_0_impl_instance: Constant_float_8_23_sinnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);

   Delay5No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => Delay5No8_out);

   Delay5No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => Delay5No9_out);

   Delay5No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => Delay5No19_out);

   Delay7No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => Delay7No_out);

   Delay7No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => Delay7No1_out);

   Delay3No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => Delay3No46_out);

   Delay4No12_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => Delay4No12_out);

   Delay4No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => Delay4No13_out);

   Delay3No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => Delay3No56_out);

   Delay3No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => Delay3No57_out);

   Delay3No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => Delay3No66_out);

   Delay3No67_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => Delay3No67_out);

   Delay5No26_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => Delay5No26_out);

   Delay5No27_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => Delay5No27_out);

   Delay3No68_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => Delay3No68_out);

   Delay5No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => Delay5No28_out);

   Delay5No29_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => Delay5No29_out);

   Delay4No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => Delay4No22_out);

   Delay4No23_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => Delay4No23_out);

   Delay3No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => Delay3No84_out);

   Delay3No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => Delay3No86_out);

   Delay3No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => Delay3No87_out);

   Delay5No30_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => Delay5No30_out);

   Delay5No31_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => Delay5No31_out);

   Delay5No32_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => Delay5No32_out);

   Delay5No33_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => Delay5No33_out);

   Delay5No34_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => Delay5No34_out);

   Delay5No35_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => Delay5No35_out);

   Delay6No6_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => Delay6No6_out);

   Delay6No7_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => Delay6No7_out);

   Delay5No36_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => Delay5No36_out);

   Delay5No37_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => Delay5No37_out);

   Delay4No32_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => Delay4No32_out);

   Delay4No33_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => Delay4No33_out);

   Delay15No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => Delay15No4_out);

   Delay15No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => Delay15No5_out);

   Delay6No8_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => Delay6No8_out);

   Delay6No9_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => Delay6No9_out);

   Delay5No41_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => Delay5No41_out);

   Delay6No10_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => Delay6No10_out);

   Delay6No11_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => Delay6No11_out);

   Delay16No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => Delay16No8_out);

   Delay16No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => Delay16No9_out);

   Delay5No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg263_out,
                 Y => Delay5No42_out);

   Delay5No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => Delay5No43_out);

   Delay5No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => Delay5No44_out);

   Delay5No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => Delay5No47_out);

   Delay5No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => Delay5No48_out);

   Delay5No49_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => Delay5No49_out);

   Delay7No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => Delay7No10_out);

   Delay7No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => Delay7No11_out);

   MUX_y0_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y0_re_0_0_LUT_out);

   MUX_y0_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y0_im_0_0_LUT_out);

   MUX_y1_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y1_re_0_0_LUT_out);

   MUX_y1_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y1_im_0_0_LUT_out);

   MUX_y2_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y2_re_0_0_LUT_out);

   MUX_y2_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y2_im_0_0_LUT_out);

   MUX_y3_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y3_re_0_0_LUT_out);

   MUX_y3_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y3_im_0_0_LUT_out);

   MUX_y4_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y4_re_0_0_LUT_out);

   MUX_y4_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y4_im_0_0_LUT_out);

   MUX_y5_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y5_re_0_0_LUT_out);

   MUX_y5_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y5_im_0_0_LUT_out);

   MUX_y6_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y6_re_0_0_LUT_out);

   MUX_y6_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y6_im_0_0_LUT_out);

   MUX_y7_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y7_re_0_0_LUT_out);

   MUX_y7_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y7_im_0_0_LUT_out);

   MUX_y8_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y8_re_0_0_LUT_out);

   MUX_y8_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y8_im_0_0_LUT_out);

   MUX_y9_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y9_re_0_0_LUT_out);

   MUX_y9_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y9_im_0_0_LUT_out);

   MUX_y10_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y10_re_0_0_LUT_out);

   MUX_y10_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y10_im_0_0_LUT_out);

   MUX_y11_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y11_re_0_0_LUT_out);

   MUX_y11_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y11_im_0_0_LUT_out);

   MUX_y12_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y12_re_0_0_LUT_out);

   MUX_y12_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y12_im_0_0_LUT_out);

   MUX_y13_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y13_re_0_0_LUT_out);

   MUX_y13_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y13_im_0_0_LUT_out);

   MUX_y14_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y14_re_0_0_LUT_out);

   MUX_y14_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y14_im_0_0_LUT_out);

   MUX_y15_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y15_re_0_0_LUT_out);

   MUX_y15_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_y15_im_0_0_LUT_out);

   MUX_Product331_1_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product331_1_impl_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_Product331_1_impl_0_LUT_out);

   MUX_Product331_1_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product331_1_impl_1_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount71_out,
                 Output => MUX_Product331_1_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_re_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_im_0_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_re_0_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_im_0_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_re_0_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_im_0_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_re_0_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_im_0_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_re_0_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_im_0_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_re_0_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_im_0_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_re_0_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_im_0_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_re_0_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_im_0_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_re_0_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_im_0_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_re_0_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_im_0_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_re_0_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_im_0_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_re_0_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_im_0_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_re_0_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_im_0_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_re_0_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_im_0_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_re_0_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_im_0_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_re_0_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_im_0_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_0_impl_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_1_impl_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_0_impl_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_1_impl_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_0_impl_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_1_impl_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_0_impl_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_1_impl_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add16_0_impl_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add16_1_impl_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_0_impl_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_1_impl_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_0_impl_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_1_impl_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add117_0_impl_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add117_1_impl_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add120_0_impl_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add120_1_impl_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add36_0_impl_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add36_1_impl_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add127_0_impl_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add127_1_impl_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add38_0_impl_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add38_1_impl_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add128_0_impl_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add128_1_impl_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add129_0_impl_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add129_1_impl_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add40_0_impl_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add40_1_impl_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add130_0_impl_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add130_1_impl_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_0_impl_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_1_impl_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_0_impl_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_1_impl_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_0_impl_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_1_impl_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_0_impl_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_1_impl_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_0_impl_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_1_impl_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_0_impl_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_1_impl_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_0_impl_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_1_impl_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_0_impl_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_1_impl_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product13_0_impl_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product13_1_impl_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_0_impl_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_1_impl_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_0_impl_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_1_impl_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_0_impl_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_1_impl_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product25_0_impl_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product25_1_impl_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product35_0_impl_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product35_1_impl_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract6_0_impl_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract6_1_impl_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product9_0_impl_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product9_1_impl_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product16_0_impl_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product16_1_impl_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_0_impl_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_1_impl_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product36_0_impl_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product36_1_impl_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract7_0_impl_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract7_1_impl_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_0_impl_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_1_impl_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_0_impl_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_1_impl_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_0_impl_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_1_impl_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_0_impl_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_1_impl_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_0_impl_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_1_impl_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract23_0_impl_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract23_1_impl_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product124_0_impl_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product124_1_impl_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product323_0_impl_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product323_1_impl_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product324_0_impl_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product324_1_impl_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product325_1_impl_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_0_impl_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product226_0_impl_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product226_1_impl_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product130_1_impl_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product329_0_impl_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product329_1_impl_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract30_0_impl_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract30_1_impl_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg332_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg334_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product132_0_impl_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product132_1_impl_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product331_0_impl_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product331_1_impl_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract42_0_impl_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg341_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract42_1_impl_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg346_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract44_0_impl_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract44_1_impl_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract45_0_impl_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg359_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg360_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract45_1_impl_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg362_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract46_0_impl_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract46_1_impl_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg369_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract57_0_impl_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg372_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract57_1_impl_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg377_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract117_0_impl_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg380_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract117_1_impl_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract61_0_impl_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract61_1_impl_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg388_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract121_0_impl_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract121_1_impl_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant2_0_impl_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg396_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => SharedReg400_out);

   SharedReg401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => SharedReg401_out);

   SharedReg402_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg401_out,
                 Y => SharedReg402_out);

   SharedReg403_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg402_out,
                 Y => SharedReg403_out);

   SharedReg404_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg403_out,
                 Y => SharedReg404_out);

   SharedReg405_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant11_0_impl_out,
                 Y => SharedReg405_out);

   SharedReg406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg405_out,
                 Y => SharedReg406_out);

   SharedReg407_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg406_out,
                 Y => SharedReg407_out);

   SharedReg408_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg407_out,
                 Y => SharedReg408_out);

   SharedReg409_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => SharedReg409_out);

   SharedReg410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg409_out,
                 Y => SharedReg410_out);

   SharedReg411_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg410_out,
                 Y => SharedReg411_out);

   SharedReg412_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg411_out,
                 Y => SharedReg412_out);

   SharedReg413_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg412_out,
                 Y => SharedReg413_out);

   SharedReg414_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg413_out,
                 Y => SharedReg414_out);

   SharedReg415_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg414_out,
                 Y => SharedReg415_out);

   SharedReg416_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg415_out,
                 Y => SharedReg416_out);

   SharedReg417_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg416_out,
                 Y => SharedReg417_out);

   SharedReg418_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant4_0_impl_out,
                 Y => SharedReg418_out);

   SharedReg419_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => SharedReg419_out);

   SharedReg420_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant13_0_impl_out,
                 Y => SharedReg420_out);

   SharedReg421_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => SharedReg421_out);

   SharedReg422_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant5_0_impl_out,
                 Y => SharedReg422_out);

   SharedReg423_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant14_0_impl_out,
                 Y => SharedReg423_out);

   SharedReg424_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant6_0_impl_out,
                 Y => SharedReg424_out);

   SharedReg425_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg424_out,
                 Y => SharedReg425_out);

   SharedReg426_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg425_out,
                 Y => SharedReg426_out);

   SharedReg427_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg426_out,
                 Y => SharedReg427_out);

   SharedReg428_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant15_0_impl_out,
                 Y => SharedReg428_out);

   SharedReg429_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => SharedReg429_out);

   SharedReg430_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg429_out,
                 Y => SharedReg430_out);

   SharedReg431_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg430_out,
                 Y => SharedReg431_out);

   SharedReg432_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant7_0_impl_out,
                 Y => SharedReg432_out);

   SharedReg433_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant16_0_impl_out,
                 Y => SharedReg433_out);

   SharedReg434_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant8_0_impl_out,
                 Y => SharedReg434_out);

   SharedReg435_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg434_out,
                 Y => SharedReg435_out);

   SharedReg436_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg435_out,
                 Y => SharedReg436_out);

   SharedReg437_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg436_out,
                 Y => SharedReg437_out);

   SharedReg438_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg437_out,
                 Y => SharedReg438_out);

   SharedReg439_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant17_0_impl_out,
                 Y => SharedReg439_out);

   SharedReg440_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => SharedReg440_out);

   SharedReg441_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg440_out,
                 Y => SharedReg441_out);

   SharedReg442_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg441_out,
                 Y => SharedReg442_out);

   SharedReg443_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => SharedReg443_out);

   SharedReg444_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant9_0_impl_out,
                 Y => SharedReg444_out);

   SharedReg445_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg444_out,
                 Y => SharedReg445_out);

   SharedReg446_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant18_0_impl_out,
                 Y => SharedReg446_out);

   SharedReg447_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg446_out,
                 Y => SharedReg447_out);

   SharedReg448_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg448_out);

   SharedReg449_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg449_out);
end architecture;

