--------------------------------------------------------------------------------
--                         ModuloCounter_28_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_28_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of ModuloCounter_28_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(4 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 27 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid175455_RightShifter
--                 (RightShifter_24_by_max_26_F250_uid175457)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid175455_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid175455_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_f250_uid175460
--                  (IntAdderAlternative_27_f250_uid175464)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid175460 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid175460 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--               LZCShifter_28_to_28_counting_32_F250_uid175467
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid175467 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid175467 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_f250_uid175470
--                   (IntAdderClassical_34_f250_uid175472)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid175470 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid175470 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                            FPAdd_8_23_uid175455
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid175455 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid175455 is
   component FPAdd_8_23_uid175455_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid175460 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid175467 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid175470 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid175455_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid175460  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid175467  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid175470  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid175455 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid175455  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_28_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_28_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(4 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_28_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00000",
         iS_1 when "00001",
         iS_2 when "00010",
         iS_3 when "00011",
         iS_4 when "00100",
         iS_5 when "00101",
         iS_6 when "00110",
         iS_7 when "00111",
         iS_8 when "01000",
         iS_9 when "01001",
         iS_10 when "01010",
         iS_11 when "01011",
         iS_12 when "01100",
         iS_13 when "01101",
         iS_14 when "01110",
         iS_15 when "01111",
         iS_16 when "10000",
         iS_17 when "10001",
         iS_18 when "10010",
         iS_19 when "10011",
         iS_20 when "10100",
         iS_21 when "10101",
         iS_22 when "10110",
         iS_23 when "10111",
         iS_24 when "11000",
         iS_25 when "11001",
         iS_26 when "11010",
         iS_27 when "11011",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid175588
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid175588 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid175588 is
signal XX_m175589 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m175589 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m175589 <= X ;
   YY_m175589 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_33_f500_uid175592
--                   (IntAdderClassical_33_f500_uid175594)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid175592 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid175592 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid175588 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid175592 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid175588  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
   RoundingAdder: IntAdder_33_f500_uid175592  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound   ,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid175631_RightShifter
--                 (RightShifter_24_by_max_26_F250_uid175633)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid175631_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid175631_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_f250_uid175636
--                  (IntAdderAlternative_27_f250_uid175640)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid175636 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid175636 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--               LZCShifter_28_to_28_counting_32_F250_uid175643
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid175643 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid175643 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_f250_uid175646
--                   (IntAdderClassical_34_f250_uid175648)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid175646 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid175646 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                            FPAdd_8_23_uid175631
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid175631 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid175631 is
   component FPAdd_8_23_uid175631_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid175636 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid175643 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid175646 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid175631_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid175636  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid175643  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid175646  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid175631 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid175631  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_26_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_26_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(4 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_26_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00000",
         iS_1 when "00001",
         iS_2 when "00010",
         iS_3 when "00011",
         iS_4 when "00100",
         iS_5 when "00101",
         iS_6 when "00110",
         iS_7 when "00111",
         iS_8 when "01000",
         iS_9 when "01001",
         iS_10 when "01010",
         iS_11 when "01011",
         iS_12 when "01100",
         iS_13 when "01101",
         iS_14 when "01110",
         iS_15 when "01111",
         iS_16 when "10000",
         iS_17 when "10001",
         iS_18 when "10010",
         iS_19 when "10011",
         iS_20 when "10100",
         iS_21 when "10101",
         iS_22 when "10110",
         iS_23 when "10111",
         iS_24 when "11000",
         iS_25 when "11001",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_0_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 23 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      Y <= s22;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 22 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      Y <= s21;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      Y <= s16;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      Y <= s17;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 25 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      Y <= s24;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 30 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      Y <= s29;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 29 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      Y <= s28;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 28 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      Y <= s27;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 27 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      Y <= s26;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 24 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      Y <= s23;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      Y <= s15;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product7_impl_0_LUT_wIn_5_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product7_impl_0_LUT_wIn_5_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product7_impl_0_LUT_wIn_5_wOut_5 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "00110" when "00000",
      "01001" when "00001",
      "01010" when "00010",
      "01011" when "00011",
      "00111" when "00100",
      "00000" when "00101",
      "01110" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "10111" when "01001",
      "10100" when "01010",
      "10101" when "01011",
      "11001" when "01100",
      "10011" when "01101",
      "10110" when "01110",
      "00010" when "01111",
      "00001" when "10000",
      "00101" when "10001",
      "11000" when "10010",
      "01101" when "10011",
      "10000" when "10100",
      "01111" when "10101",
      "10001" when "10110",
      "01100" when "10111",
      "00011" when "11000",
      "10010" when "11001",
      "01000" when "11010",
      "00100" when "11011",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product7_impl_0_LUT_wIn_5_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product7_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product7_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product7_impl_0_LUT_wIn_5_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_Product7_impl_0_LUT_wIn_5_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product7_impl_1_LUT_wIn_5_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product7_impl_1_LUT_wIn_5_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product7_impl_1_LUT_wIn_5_wOut_5 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "01000" when "00000",
      "10100" when "00001",
      "10101" when "00010",
      "01010" when "00011",
      "01001" when "00100",
      "10110" when "00101",
      "00001" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00101" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00111" when "01100",
      "10010" when "01101",
      "00100" when "01110",
      "10111" when "01111",
      "11000" when "10000",
      "10011" when "10001",
      "00110" when "10010",
      "01101" when "10011",
      "01110" when "10100",
      "10000" when "10101",
      "01111" when "10110",
      "01100" when "10111",
      "11001" when "11000",
      "10001" when "11001",
      "00000" when "11010",
      "01011" when "11011",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product7_impl_1_LUT_wIn_5_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product7_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product7_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product7_impl_1_LUT_wIn_5_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_Product7_impl_1_LUT_wIn_5_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product220_impl_0_LUT_wIn_5_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product220_impl_0_LUT_wIn_5_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product220_impl_0_LUT_wIn_5_wOut_5 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "01001" when "00000",
      "01010" when "00001",
      "01011" when "00010",
      "01100" when "00011",
      "00100" when "00100",
      "01101" when "00101",
      "11000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00000" when "01010",
      "10111" when "01011",
      "00011" when "01100",
      "10011" when "01101",
      "00001" when "01110",
      "01110" when "01111",
      "10101" when "10000",
      "10110" when "10001",
      "11001" when "10010",
      "01111" when "10011",
      "00111" when "10100",
      "10001" when "10101",
      "10000" when "10110",
      "00110" when "10111",
      "10100" when "11000",
      "01000" when "11001",
      "10010" when "11010",
      "00101" when "11011",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product220_impl_0_LUT_wIn_5_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product220_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product220_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product220_impl_0_LUT_wIn_5_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_Product220_impl_0_LUT_wIn_5_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product220_impl_1_LUT_wIn_5_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product220_impl_1_LUT_wIn_5_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product220_impl_1_LUT_wIn_5_wOut_5 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "00111" when "00000",
      "10000" when "00001",
      "10001" when "00010",
      "01001" when "00011",
      "10010" when "00100",
      "01000" when "00101",
      "00101" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "11000" when "01001",
      "10110" when "01010",
      "00100" when "01011",
      "11001" when "01100",
      "01110" when "01101",
      "10111" when "01110",
      "01010" when "01111",
      "00010" when "10000",
      "00011" when "10001",
      "00110" when "10010",
      "01011" when "10011",
      "10100" when "10100",
      "00001" when "10101",
      "01100" when "10110",
      "10011" when "10111",
      "01101" when "11000",
      "10101" when "11001",
      "00000" when "11010",
      "01111" when "11011",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product220_impl_1_LUT_wIn_5_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product220_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product220_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product220_impl_1_LUT_wIn_5_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_Product220_impl_1_LUT_wIn_5_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 43 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      Y <= s42;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 56 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      Y <= s55;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 58 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      Y <= s57;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 57 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      Y <= s56;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 54 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      Y <= s53;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 36 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      Y <= s35;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 33 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      Y <= s32;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 31 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      Y <= s30;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 32 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      Y <= s31;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 55 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      Y <= s54;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 60 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      Y <= s59;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 34 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      Y <= s33;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_79_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 79 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_79_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_79_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      Y <= s78;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_77_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 77 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_77_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_77_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      Y <= s76;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 78 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      Y <= s77;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 104 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      Y <= s103;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 99 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      Y <= s98;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 76 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      Y <= s75;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_100_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 100 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_100_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_100_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      Y <= s99;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 69 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      Y <= s68;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 53 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      Y <= s52;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 81 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      Y <= s80;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          x0_re : in std_logic_vector(31 downto 0);
          x0_im : in std_logic_vector(31 downto 0);
          x1_re : in std_logic_vector(31 downto 0);
          x1_im : in std_logic_vector(31 downto 0);
          x2_re : in std_logic_vector(31 downto 0);
          x2_im : in std_logic_vector(31 downto 0);
          x3_re : in std_logic_vector(31 downto 0);
          x3_im : in std_logic_vector(31 downto 0);
          x4_re : in std_logic_vector(31 downto 0);
          x4_im : in std_logic_vector(31 downto 0);
          x5_re : in std_logic_vector(31 downto 0);
          x5_im : in std_logic_vector(31 downto 0);
          x6_re : in std_logic_vector(31 downto 0);
          x6_im : in std_logic_vector(31 downto 0);
          x7_re : in std_logic_vector(31 downto 0);
          x7_im : in std_logic_vector(31 downto 0);
          x8_re : in std_logic_vector(31 downto 0);
          x8_im : in std_logic_vector(31 downto 0);
          x9_re : in std_logic_vector(31 downto 0);
          x9_im : in std_logic_vector(31 downto 0);
          x10_re : in std_logic_vector(31 downto 0);
          x10_im : in std_logic_vector(31 downto 0);
          x11_re : in std_logic_vector(31 downto 0);
          x11_im : in std_logic_vector(31 downto 0);
          x12_re : in std_logic_vector(31 downto 0);
          x12_im : in std_logic_vector(31 downto 0);
          x13_re : in std_logic_vector(31 downto 0);
          x13_im : in std_logic_vector(31 downto 0);
          x14_re : in std_logic_vector(31 downto 0);
          x14_im : in std_logic_vector(31 downto 0);
          x15_re : in std_logic_vector(31 downto 0);
          x15_im : in std_logic_vector(31 downto 0);
          y0_re : out std_logic_vector(31 downto 0);
          y0_im : out std_logic_vector(31 downto 0);
          y1_re : out std_logic_vector(31 downto 0);
          y1_im : out std_logic_vector(31 downto 0);
          y2_re : out std_logic_vector(31 downto 0);
          y2_im : out std_logic_vector(31 downto 0);
          y3_re : out std_logic_vector(31 downto 0);
          y3_im : out std_logic_vector(31 downto 0);
          y4_re : out std_logic_vector(31 downto 0);
          y4_im : out std_logic_vector(31 downto 0);
          y5_re : out std_logic_vector(31 downto 0);
          y5_im : out std_logic_vector(31 downto 0);
          y6_re : out std_logic_vector(31 downto 0);
          y6_im : out std_logic_vector(31 downto 0);
          y7_re : out std_logic_vector(31 downto 0);
          y7_im : out std_logic_vector(31 downto 0);
          y8_re : out std_logic_vector(31 downto 0);
          y8_im : out std_logic_vector(31 downto 0);
          y9_re : out std_logic_vector(31 downto 0);
          y9_im : out std_logic_vector(31 downto 0);
          y10_re : out std_logic_vector(31 downto 0);
          y10_im : out std_logic_vector(31 downto 0);
          y11_re : out std_logic_vector(31 downto 0);
          y11_im : out std_logic_vector(31 downto 0);
          y12_re : out std_logic_vector(31 downto 0);
          y12_im : out std_logic_vector(31 downto 0);
          y13_re : out std_logic_vector(31 downto 0);
          y13_im : out std_logic_vector(31 downto 0);
          y14_re : out std_logic_vector(31 downto 0);
          y14_im : out std_logic_vector(31 downto 0);
          y15_re : out std_logic_vector(31 downto 0);
          y15_im : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_28_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(4 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_28_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(4 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_26_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(4 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product7_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product7_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product220_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product220_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_79_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_77_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_100_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount281_out : std_logic_vector(4 downto 0) := (others => '0');
signal x0_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add120_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add120_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add120_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product13_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract17_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract17_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract17_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract20_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product220_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product220_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product220_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant11_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant12_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant13_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant14_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant15_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant16_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant17_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant9_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant18_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant10_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant19_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant20_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant110_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant21_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant111_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant22_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant112_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant23_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant113_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant24_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant114_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant25_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant115_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant26_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant116_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant27_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant117_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant28_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant118_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant29_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant119_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant30_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant120_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant31_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant121_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant32_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant122_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant33_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant123_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant34_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant124_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant35_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant125_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant36_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant126_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant37_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant127_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant38_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant128_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant39_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant129_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant40_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant130_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant41_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant131_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant42_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant132_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant43_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant133_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant44_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant134_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant45_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant135_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant46_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant136_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant47_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant137_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant48_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant138_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant49_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant139_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant50_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant140_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant51_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant141_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant52_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant142_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant53_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant143_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant54_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant144_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant55_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant145_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant56_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant146_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant57_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant147_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay28No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay29No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay33No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay33No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay30No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay28No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay24No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay29No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay29No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay30No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay31No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay34No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay34No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay60No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay60No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay35No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay57No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay57No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay39No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay54No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay54No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay54No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay55No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay63No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay62No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay57No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay57No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay63No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay55No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay35No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay35No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay105No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay105No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay34No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay69No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay82No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay69No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay38No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay42No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay42No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product7_impl_0_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product7_impl_1_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product220_impl_0_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product220_impl_1_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x0_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y1_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y1_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y2_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y2_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y3_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y3_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y4_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y4_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y5_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y5_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y6_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y6_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y7_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y7_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y8_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y8_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y9_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y9_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y10_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y10_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y11_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y11_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y12_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y12_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y13_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y13_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y14_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y14_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y15_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y15_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No32_out_to_Add2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Add2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No1_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No1_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay30No1_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No3_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No4_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No2_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No1_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No1_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No6_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Add7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Add7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Add9_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Add9_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No1_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay29No15_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Add120_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Add120_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No3_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay33No_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No7_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay29No2_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Product4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Product4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay57No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay34No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay35No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No17_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No5_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No5_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No2_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay54No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay55No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No14_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Product21_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Product21_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay57No1_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay63No_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No19_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No9_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No6_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No3_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay34No1_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No1_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay33No1_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Product13_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Product13_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay62No_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay69No2_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No5_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No10_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay105No_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No3_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No1_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay63No1_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No20_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No2_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No7_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Product23_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Product23_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No1_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay35No2_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay39No_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No2_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No6_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No1_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No2_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No6_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No1_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay54No3_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay55No6_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay28No2_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay105No1_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Product33_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Product33_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No2_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No1_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No1_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay69No5_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No3_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No2_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No4_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay54No4_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay35No1_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No7_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Subtract4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Subtract4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No1_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay28No3_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No3_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No5_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Product7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Product7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay60No_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay57No3_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay34No4_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No6_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No3_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay42No_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No10_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay30No2_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No5_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Subtract17_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Subtract17_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No2_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay24No3_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No7_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay29No17_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Subtract20_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Subtract20_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No3_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No2_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No7_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Product220_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Product220_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay57No4_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No3_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No1_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay82No_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No6_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No8_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No11_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay31No_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay60No1_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No4_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay38No_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay42No1_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount281_instance: ModuloCounter_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount281_out);
x0_re_IEEE <= x0_re;
   x0_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_re_out,
                 X => x0_re_IEEE);
x0_im_IEEE <= x0_im;
   x0_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_im_out,
                 X => x0_im_IEEE);
x1_re_IEEE <= x1_re;
   x1_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_re_out,
                 X => x1_re_IEEE);
x1_im_IEEE <= x1_im;
   x1_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_im_out,
                 X => x1_im_IEEE);
x2_re_IEEE <= x2_re;
   x2_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_re_out,
                 X => x2_re_IEEE);
x2_im_IEEE <= x2_im;
   x2_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_im_out,
                 X => x2_im_IEEE);
x3_re_IEEE <= x3_re;
   x3_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_re_out,
                 X => x3_re_IEEE);
x3_im_IEEE <= x3_im;
   x3_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_im_out,
                 X => x3_im_IEEE);
x4_re_IEEE <= x4_re;
   x4_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_re_out,
                 X => x4_re_IEEE);
x4_im_IEEE <= x4_im;
   x4_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_im_out,
                 X => x4_im_IEEE);
x5_re_IEEE <= x5_re;
   x5_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_re_out,
                 X => x5_re_IEEE);
x5_im_IEEE <= x5_im;
   x5_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_im_out,
                 X => x5_im_IEEE);
x6_re_IEEE <= x6_re;
   x6_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_re_out,
                 X => x6_re_IEEE);
x6_im_IEEE <= x6_im;
   x6_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_im_out,
                 X => x6_im_IEEE);
x7_re_IEEE <= x7_re;
   x7_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_re_out,
                 X => x7_re_IEEE);
x7_im_IEEE <= x7_im;
   x7_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_im_out,
                 X => x7_im_IEEE);
x8_re_IEEE <= x8_re;
   x8_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_re_out,
                 X => x8_re_IEEE);
x8_im_IEEE <= x8_im;
   x8_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_im_out,
                 X => x8_im_IEEE);
x9_re_IEEE <= x9_re;
   x9_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_re_out,
                 X => x9_re_IEEE);
x9_im_IEEE <= x9_im;
   x9_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_im_out,
                 X => x9_im_IEEE);
x10_re_IEEE <= x10_re;
   x10_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_re_out,
                 X => x10_re_IEEE);
x10_im_IEEE <= x10_im;
   x10_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_im_out,
                 X => x10_im_IEEE);
x11_re_IEEE <= x11_re;
   x11_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_re_out,
                 X => x11_re_IEEE);
x11_im_IEEE <= x11_im;
   x11_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_im_out,
                 X => x11_im_IEEE);
x12_re_IEEE <= x12_re;
   x12_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_re_out,
                 X => x12_re_IEEE);
x12_im_IEEE <= x12_im;
   x12_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_im_out,
                 X => x12_im_IEEE);
x13_re_IEEE <= x13_re;
   x13_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_re_out,
                 X => x13_re_IEEE);
x13_im_IEEE <= x13_im;
   x13_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_im_out,
                 X => x13_im_IEEE);
x14_re_IEEE <= x14_re;
   x14_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_re_out,
                 X => x14_re_IEEE);
x14_im_IEEE <= x14_im;
   x14_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_im_out,
                 X => x14_im_IEEE);
x15_re_IEEE <= x15_re;
   x15_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_re_out,
                 X => x15_re_IEEE);
x15_im_IEEE <= x15_im;
   x15_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_im_out,
                 X => x15_im_IEEE);
   y0_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_re_IEEE,
                 X => Delay1No_out);
y0_re <= y0_re_IEEE;

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => Delay1No_out);
   y0_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_im_IEEE,
                 X => Delay1No1_out);
y0_im <= y0_im_IEEE;

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => Delay1No1_out);
   y1_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_re_IEEE,
                 X => Delay1No2_out);
y1_re <= y1_re_IEEE;

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => Delay1No2_out);
   y1_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_im_IEEE,
                 X => Delay1No3_out);
y1_im <= y1_im_IEEE;

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => Delay1No3_out);
   y2_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_re_IEEE,
                 X => Delay1No4_out);
y2_re <= y2_re_IEEE;

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => Delay1No4_out);
   y2_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_im_IEEE,
                 X => Delay1No5_out);
y2_im <= y2_im_IEEE;

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => Delay1No5_out);
   y3_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_re_IEEE,
                 X => Delay1No6_out);
y3_re <= y3_re_IEEE;

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => Delay1No6_out);
   y3_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_im_IEEE,
                 X => Delay1No7_out);
y3_im <= y3_im_IEEE;

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => Delay1No7_out);
   y4_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_re_IEEE,
                 X => Delay1No8_out);
y4_re <= y4_re_IEEE;

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => Delay1No8_out);
   y4_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_im_IEEE,
                 X => Delay1No9_out);
y4_im <= y4_im_IEEE;

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => Delay1No9_out);
   y5_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_re_IEEE,
                 X => Delay1No10_out);
y5_re <= y5_re_IEEE;

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => Delay1No10_out);
   y5_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_im_IEEE,
                 X => Delay1No11_out);
y5_im <= y5_im_IEEE;

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => Delay1No11_out);
   y6_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_re_IEEE,
                 X => Delay1No12_out);
y6_re <= y6_re_IEEE;

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => Delay1No12_out);
   y6_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_im_IEEE,
                 X => Delay1No13_out);
y6_im <= y6_im_IEEE;

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => Delay1No13_out);
   y7_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_re_IEEE,
                 X => Delay1No14_out);
y7_re <= y7_re_IEEE;

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => Delay1No14_out);
   y7_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_im_IEEE,
                 X => Delay1No15_out);
y7_im <= y7_im_IEEE;

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => Delay1No15_out);
   y8_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_re_IEEE,
                 X => Delay1No16_out);
y8_re <= y8_re_IEEE;

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => Delay1No16_out);
   y8_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_im_IEEE,
                 X => Delay1No17_out);
y8_im <= y8_im_IEEE;

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => Delay1No17_out);
   y9_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_re_IEEE,
                 X => Delay1No18_out);
y9_re <= y9_re_IEEE;

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => Delay1No18_out);
   y9_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_im_IEEE,
                 X => Delay1No19_out);
y9_im <= y9_im_IEEE;

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => Delay1No19_out);
   y10_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_re_IEEE,
                 X => Delay1No20_out);
y10_re <= y10_re_IEEE;

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => Delay1No20_out);
   y10_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_im_IEEE,
                 X => Delay1No21_out);
y10_im <= y10_im_IEEE;

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => Delay1No21_out);
   y11_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_re_IEEE,
                 X => Delay1No22_out);
y11_re <= y11_re_IEEE;

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => Delay1No22_out);
   y11_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_im_IEEE,
                 X => Delay1No23_out);
y11_im <= y11_im_IEEE;

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => Delay1No23_out);
   y12_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_re_IEEE,
                 X => Delay1No24_out);
y12_re <= y12_re_IEEE;

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => Delay1No24_out);
   y12_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_im_IEEE,
                 X => Delay1No25_out);
y12_im <= y12_im_IEEE;

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => Delay1No25_out);
   y13_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_re_IEEE,
                 X => Delay1No26_out);
y13_re <= y13_re_IEEE;

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => Delay1No26_out);
   y13_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_im_IEEE,
                 X => Delay1No27_out);
y13_im <= y13_im_IEEE;

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => Delay1No27_out);
   y14_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_re_IEEE,
                 X => Delay1No28_out);
y14_re <= y14_re_IEEE;

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => Delay1No28_out);
   y14_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_im_IEEE,
                 X => Delay1No29_out);
y14_im <= y14_im_IEEE;

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => Delay1No29_out);
   y15_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_re_IEEE,
                 X => Delay1No30_out);
y15_re <= y15_re_IEEE;

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => Delay1No30_out);
   y15_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_im_IEEE,
                 X => Delay1No31_out);
y15_im <= y15_im_IEEE;

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Add2_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Add2_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Add2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_impl_out,
                 X => Delay1No32_out_to_Add2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Add2_impl_parent_implementedSystem_port_1_cast);

SharedReg48_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg48_out;
SharedReg4_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg4_out;
SharedReg128_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg128_out;
SharedReg117_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg117_out;
SharedReg5_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg5_out;
SharedReg65_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg65_out;
Delay6No1_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_7_cast <= Delay6No1_out;
Delay7No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_8_cast <= Delay7No_out;
Delay8No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_9_cast <= Delay8No_out;
Delay9No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_10_cast <= Delay9No_out;
Delay10No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_11_cast <= Delay10No_out;
SharedReg2_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg2_out;
Delay12No1_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_13_cast <= Delay12No1_out;
Delay30No1_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_14_cast <= Delay30No1_out;
SharedReg48_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg48_out;
SharedReg124_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg124_out;
SharedReg97_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg97_out;
SharedReg65_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg65_out;
SharedReg121_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg121_out;
SharedReg116_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg116_out;
SharedReg118_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg118_out;
SharedReg84_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg84_out;
SharedReg65_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg65_out;
SharedReg82_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg82_out;
SharedReg48_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg48_out;
SharedReg171_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg171_out;
SharedReg65_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg65_out;
SharedReg169_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg169_out;
   MUX_Add2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg48_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg4_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay10No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg2_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay12No1_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay30No1_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg48_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg124_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg97_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg65_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg121_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg116_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg128_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg118_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg84_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg65_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg82_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg48_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg171_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg65_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg169_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg117_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg5_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg65_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay6No1_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay7No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay8No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay9No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_impl_0_out,
                 Y => Delay1No32_out);

SharedReg69_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg69_out;
SharedReg20_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg117_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg117_out;
SharedReg165_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg165_out;
SharedReg21_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg21_out;
SharedReg82_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg82_out;
Delay6No3_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_7_cast <= Delay6No3_out;
Delay7No4_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_8_cast <= Delay7No4_out;
Delay8No2_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_9_cast <= Delay8No2_out;
Delay9No1_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_10_cast <= Delay9No1_out;
Delay10No1_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_11_cast <= Delay10No1_out;
SharedReg18_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg18_out;
Delay12No6_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_13_cast <= Delay12No6_out;
SharedReg95_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg95_out;
SharedReg81_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg81_out;
SharedReg174_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg174_out;
SharedReg132_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg132_out;
SharedReg83_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg83_out;
SharedReg117_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg117_out;
SharedReg96_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg96_out;
SharedReg166_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg166_out;
SharedReg32_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg32_out;
SharedReg82_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg82_out;
SharedReg89_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg89_out;
SharedReg82_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg82_out;
SharedReg165_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg165_out;
SharedReg87_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg87_out;
SharedReg191_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg191_out;
   MUX_Add2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay10No1_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg18_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay12No6_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg95_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg81_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg174_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg132_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg83_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg117_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg96_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg117_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg166_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg32_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg82_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg89_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg82_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg165_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg87_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg191_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg165_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg21_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg82_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay6No3_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay7No4_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay8No2_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay9No1_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Add7_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Add7_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Add7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add7_impl_out,
                 X => Delay1No34_out_to_Add7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Add7_impl_parent_implementedSystem_port_1_cast);

SharedReg65_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg65_out;
SharedReg93_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg93_out;
SharedReg153_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg153_out;
SharedReg82_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg82_out;
SharedReg117_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg117_out;
SharedReg9_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg9_out;
SharedReg123_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg123_out;
SharedReg48_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg48_out;
SharedReg200_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg200_out;
SharedReg145_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg145_out;
SharedReg135_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg135_out;
SharedReg7_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg7_out;
SharedReg14_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg14_out;
SharedReg120_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg120_out;
SharedReg169_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg169_out;
SharedReg117_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg117_out;
SharedReg96_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg96_out;
SharedReg108_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg108_out;
SharedReg88_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg88_out;
SharedReg141_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg141_out;
SharedReg85_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg85_out;
SharedReg187_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg187_out;
SharedReg96_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg96_out;
SharedReg108_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg108_out;
SharedReg117_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg117_out;
SharedReg65_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg65_out;
SharedReg165_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg165_out;
SharedReg82_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg82_out;
   MUX_Add7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg65_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg93_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg135_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg7_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg14_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg120_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg169_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg117_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg96_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg108_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg88_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg141_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg153_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg85_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg187_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg96_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg108_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg117_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg65_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg165_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg82_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg82_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg117_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg9_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg123_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg48_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg200_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg145_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add7_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add7_impl_0_out,
                 Y => Delay1No34_out);

SharedReg82_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg82_out;
SharedReg72_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg72_out;
SharedReg96_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg96_out;
SharedReg90_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg90_out;
SharedReg165_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg165_out;
SharedReg25_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg117_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg117_out;
SharedReg65_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg65_out;
SharedReg117_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg117_out;
SharedReg223_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg223_out;
SharedReg147_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg147_out;
SharedReg23_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg23_out;
SharedReg30_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg30_out;
SharedReg117_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg117_out;
SharedReg128_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg128_out;
SharedReg204_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg204_out;
SharedReg108_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg108_out;
SharedReg130_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg130_out;
SharedReg82_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg82_out;
SharedReg148_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg148_out;
SharedReg87_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg87_out;
SharedReg117_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg117_out;
SharedReg102_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg102_out;
SharedReg159_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg159_out;
SharedReg165_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg165_out;
SharedReg82_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg82_out;
SharedReg120_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg120_out;
SharedReg53_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg53_out;
   MUX_Add7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg82_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg147_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg23_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg30_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg117_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg128_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg204_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg108_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg130_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg82_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg148_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg96_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg87_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg117_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg102_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg159_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg165_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg82_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg120_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg53_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg90_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg165_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg25_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg117_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg65_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg117_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg223_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add7_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add7_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Add9_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Add9_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Add9_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_impl_out,
                 X => Delay1No36_out_to_Add9_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Add9_impl_parent_implementedSystem_port_1_cast);

SharedReg130_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_1_cast <= SharedReg130_out;
SharedReg129_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_2_cast <= SharedReg129_out;
SharedReg114_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_3_cast <= SharedReg114_out;
SharedReg106_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_4_cast <= SharedReg106_out;
SharedReg193_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_5_cast <= SharedReg193_out;
SharedReg11_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_6_cast <= SharedReg11_out;
SharedReg173_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_7_cast <= SharedReg173_out;
SharedReg57_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_8_cast <= SharedReg57_out;
SharedReg65_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_9_cast <= SharedReg65_out;
SharedReg141_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_10_cast <= SharedReg141_out;
SharedReg181_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_11_cast <= SharedReg181_out;
SharedReg15_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_12_cast <= SharedReg15_out;
SharedReg101_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_13_cast <= SharedReg101_out;
Delay13No_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_14_cast <= Delay13No_out;
SharedReg117_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_15_cast <= SharedReg117_out;
SharedReg48_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_16_cast <= SharedReg48_out;
SharedReg161_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_17_cast <= SharedReg161_out;
SharedReg228_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_18_cast <= SharedReg228_out;
SharedReg122_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_19_cast <= SharedReg122_out;
SharedReg142_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_20_cast <= SharedReg142_out;
SharedReg141_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_21_cast <= SharedReg141_out;
SharedReg130_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_22_cast <= SharedReg130_out;
SharedReg108_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_23_cast <= SharedReg108_out;
SharedReg141_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_24_cast <= SharedReg141_out;
SharedReg118_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_25_cast <= SharedReg118_out;
SharedReg117_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_26_cast <= SharedReg117_out;
SharedReg129_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_27_cast <= SharedReg129_out;
SharedReg48_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_28_cast <= SharedReg48_out;
   MUX_Add9_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg130_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg129_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg181_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg15_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg101_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay13No_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg117_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg48_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg161_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg228_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg122_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg142_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg114_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg141_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg130_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg108_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg141_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg118_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg117_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg129_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg48_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg106_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg193_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg11_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg173_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg57_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg65_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg141_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add9_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_impl_0_out,
                 Y => Delay1No36_out);

SharedReg141_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_1_cast <= SharedReg141_out;
SharedReg172_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_2_cast <= SharedReg172_out;
SharedReg115_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_3_cast <= SharedReg115_out;
SharedReg108_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_4_cast <= SharedReg108_out;
SharedReg210_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_5_cast <= SharedReg210_out;
SharedReg27_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_6_cast <= SharedReg27_out;
SharedReg165_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_7_cast <= SharedReg165_out;
SharedReg82_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_8_cast <= SharedReg82_out;
SharedReg82_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_9_cast <= SharedReg82_out;
SharedReg154_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_10_cast <= SharedReg154_out;
SharedReg156_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_11_cast <= SharedReg156_out;
SharedReg31_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_12_cast <= SharedReg31_out;
SharedReg108_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_13_cast <= SharedReg108_out;
Delay13No1_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_14_cast <= Delay13No1_out;
SharedReg165_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_15_cast <= SharedReg165_out;
SharedReg65_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_16_cast <= SharedReg65_out;
SharedReg130_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_17_cast <= SharedReg130_out;
Delay29No15_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_18_cast <= Delay29No15_out;
SharedReg168_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_19_cast <= SharedReg168_out;
SharedReg223_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_20_cast <= SharedReg223_out;
SharedReg154_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_21_cast <= SharedReg154_out;
SharedReg141_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_22_cast <= SharedReg141_out;
SharedReg130_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_23_cast <= SharedReg130_out;
SharedReg154_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_24_cast <= SharedReg154_out;
SharedReg202_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_25_cast <= SharedReg202_out;
SharedReg192_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_26_cast <= SharedReg192_out;
SharedReg170_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_27_cast <= SharedReg170_out;
SharedReg65_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_28_cast <= SharedReg65_out;
   MUX_Add9_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg141_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg172_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg156_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg31_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg108_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay13No1_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg165_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg65_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg130_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => Delay29No15_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg168_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg223_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg115_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg154_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg141_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg130_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg154_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg202_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg192_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg170_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg65_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg108_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg210_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg27_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg165_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg82_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg82_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg154_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add9_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Add120_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Add120_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Add120_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add120_impl_out,
                 X => Delay1No38_out_to_Add120_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Add120_impl_parent_implementedSystem_port_1_cast);

SharedReg96_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_1_cast <= SharedReg96_out;
SharedReg145_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_2_cast <= SharedReg145_out;
SharedReg224_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_3_cast <= SharedReg224_out;
SharedReg154_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_4_cast <= SharedReg154_out;
SharedReg95_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_5_cast <= SharedReg95_out;
Delay5No3_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_6_cast <= Delay5No3_out;
SharedReg98_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_7_cast <= SharedReg98_out;
SharedReg177_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_8_cast <= SharedReg177_out;
SharedReg176_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_9_cast <= SharedReg176_out;
SharedReg221_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_10_cast <= SharedReg221_out;
SharedReg152_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_11_cast <= SharedReg152_out;
SharedReg132_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_12_cast <= SharedReg132_out;
SharedReg134_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_13_cast <= SharedReg134_out;
Delay33No_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_14_cast <= Delay33No_out;
SharedReg155_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_15_cast <= SharedReg155_out;
SharedReg108_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_16_cast <= SharedReg108_out;
SharedReg229_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_17_cast <= SharedReg229_out;
SharedReg186_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_18_cast <= SharedReg186_out;
SharedReg102_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_19_cast <= SharedReg102_out;
SharedReg164_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_20_cast <= SharedReg164_out;
SharedReg184_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_21_cast <= SharedReg184_out;
SharedReg180_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_22_cast <= SharedReg180_out;
SharedReg179_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_23_cast <= SharedReg179_out;
SharedReg176_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_24_cast <= SharedReg176_out;
SharedReg32_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_25_cast <= SharedReg32_out;
SharedReg130_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_26_cast <= SharedReg130_out;
SharedReg186_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_27_cast <= SharedReg186_out;
SharedReg130_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_28_cast <= SharedReg130_out;
   MUX_Add120_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg96_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg145_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg152_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg132_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg134_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay33No_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg155_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg108_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg229_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg186_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg102_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg164_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg224_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg184_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg180_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg179_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg176_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg32_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg130_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg186_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg130_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg154_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg95_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay5No3_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg98_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg177_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg176_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg221_out_to_MUX_Add120_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add120_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add120_impl_0_out,
                 Y => Delay1No38_out);

SharedReg108_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_1_cast <= SharedReg108_out;
SharedReg108_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_2_cast <= SharedReg108_out;
SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_3_cast <= SharedReg221_out;
SharedReg176_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_4_cast <= SharedReg176_out;
SharedReg84_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_5_cast <= SharedReg84_out;
Delay5No7_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_6_cast <= Delay5No7_out;
SharedReg109_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_7_cast <= SharedReg109_out;
SharedReg222_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_8_cast <= SharedReg222_out;
SharedReg223_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_9_cast <= SharedReg223_out;
SharedReg178_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_10_cast <= SharedReg178_out;
SharedReg176_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_11_cast <= SharedReg176_out;
SharedReg144_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_12_cast <= SharedReg144_out;
SharedReg146_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_13_cast <= SharedReg146_out;
SharedReg132_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_14_cast <= SharedReg132_out;
SharedReg177_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_15_cast <= SharedReg177_out;
SharedReg131_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_16_cast <= SharedReg131_out;
SharedReg183_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_17_cast <= SharedReg183_out;
SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_18_cast <= SharedReg221_out;
Delay29No2_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_19_cast <= Delay29No2_out;
SharedReg226_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_20_cast <= SharedReg226_out;
SharedReg163_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_21_cast <= SharedReg163_out;
SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_22_cast <= SharedReg221_out;
SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_23_cast <= SharedReg221_out;
SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_24_cast <= SharedReg221_out;
SharedReg94_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_25_cast <= SharedReg94_out;
SharedReg109_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_26_cast <= SharedReg109_out;
SharedReg149_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_27_cast <= SharedReg149_out;
SharedReg141_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_28_cast <= SharedReg141_out;
   MUX_Add120_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg108_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg108_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg176_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg144_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg146_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg132_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg177_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg131_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg183_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => Delay29No2_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg226_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg163_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg221_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg94_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg109_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg149_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg141_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg176_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg84_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay5No7_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg109_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg222_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg223_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg178_out_to_MUX_Add120_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add120_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add120_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Product4_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Product4_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Product4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_impl_out,
                 X => Delay1No40_out_to_Product4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Product4_impl_parent_implementedSystem_port_1_cast);

SharedReg248_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg248_out;
Delay57No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_2_cast <= Delay57No_out;
SharedReg250_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg250_out;
Delay59No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_4_cast <= Delay59No_out;
SharedReg264_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg264_out;
SharedReg32_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg32_out;
Delay34No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_7_cast <= Delay34No_out;
Delay35No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_8_cast <= Delay35No_out;
SharedReg216_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg216_out;
SharedReg46_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg46_out;
SharedReg239_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg239_out;
Delay11No17_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_12_cast <= Delay11No17_out;
SharedReg242_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg242_out;
SharedReg310_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg310_out;
SharedReg232_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg232_out;
SharedReg235_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg235_out;
SharedReg234_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg234_out;
SharedReg188_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg188_out;
Delay18No5_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_19_cast <= Delay18No5_out;
Delay19No5_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_20_cast <= Delay19No5_out;
SharedReg292_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg292_out;
SharedReg286_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg286_out;
SharedReg32_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg32_out;
SharedReg284_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg284_out;
Delay80No2_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_25_cast <= Delay80No2_out;
SharedReg48_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg48_out;
Delay54No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_27_cast <= Delay54No_out;
Delay55No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_28_cast <= Delay55No_out;
   MUX_Product4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg248_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay57No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg239_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay11No17_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg242_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg310_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg232_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg235_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg234_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg188_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => Delay18No5_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay19No5_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg250_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg292_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg286_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg32_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg284_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => Delay80No2_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg48_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => Delay54No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => Delay55No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => Delay59No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg264_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg32_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay34No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay35No_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg216_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg46_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_impl_0_out,
                 Y => Delay1No40_out);

SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg32_out;
SharedReg65_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg65_out;
SharedReg65_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg65_out;
SharedReg84_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg84_out;
SharedReg203_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg203_out;
SharedReg267_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg267_out;
SharedReg44_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg44_out;
SharedReg215_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg215_out;
Delay36No_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_9_cast <= Delay36No_out;
Delay37No_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_10_cast <= Delay37No_out;
SharedReg206_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg206_out;
SharedReg203_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg203_out;
SharedReg203_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg203_out;
SharedReg48_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg48_out;
SharedReg33_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg33_out;
SharedReg47_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg47_out;
SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg32_out;
Delay17No14_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_18_cast <= Delay17No14_out;
SharedReg189_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg189_out;
SharedReg193_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg193_out;
SharedReg49_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg49_out;
SharedReg49_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg49_out;
SharedReg287_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg287_out;
SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg32_out;
SharedReg34_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg34_out;
SharedReg311_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg311_out;
SharedReg45_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg45_out;
SharedReg165_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg165_out;
   MUX_Product4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg65_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg206_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg203_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg203_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg48_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg33_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg47_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => Delay17No14_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg189_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg193_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg65_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg49_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg49_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg287_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg34_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg311_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg45_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg165_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg84_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg203_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg267_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg44_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg215_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay36No_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay37No_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Product21_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Product21_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Product21_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_impl_out,
                 X => Delay1No42_out_to_Product21_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Product21_impl_parent_implementedSystem_port_1_cast);

SharedReg32_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
Delay57No1_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_2_cast <= Delay57No1_out;
SharedReg262_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_3_cast <= SharedReg262_out;
SharedReg259_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_4_cast <= SharedReg259_out;
SharedReg268_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_5_cast <= SharedReg268_out;
SharedReg258_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_6_cast <= SharedReg258_out;
SharedReg218_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_7_cast <= SharedReg218_out;
Delay63No_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_8_cast <= Delay63No_out;
Delay64No_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_9_cast <= Delay64No_out;
SharedReg240_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_10_cast <= SharedReg240_out;
SharedReg276_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_11_cast <= SharedReg276_out;
Delay11No19_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_12_cast <= Delay11No19_out;
SharedReg243_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_13_cast <= SharedReg243_out;
SharedReg310_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_14_cast <= SharedReg310_out;
SharedReg233_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_15_cast <= SharedReg233_out;
SharedReg236_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_16_cast <= SharedReg236_out;
SharedReg47_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_17_cast <= SharedReg47_out;
Delay17No9_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_18_cast <= Delay17No9_out;
SharedReg246_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_19_cast <= SharedReg246_out;
Delay19No6_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_20_cast <= Delay19No6_out;
SharedReg293_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_21_cast <= SharedReg293_out;
SharedReg34_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_22_cast <= SharedReg34_out;
SharedReg56_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_23_cast <= SharedReg56_out;
SharedReg48_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_24_cast <= SharedReg48_out;
Delay80No3_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_25_cast <= Delay80No3_out;
Delay81No_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_26_cast <= Delay81No_out;
SharedReg254_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_27_cast <= SharedReg254_out;
SharedReg265_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_28_cast <= SharedReg265_out;
   MUX_Product21_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay57No1_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg276_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay11No19_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg243_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg310_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg233_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg236_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg47_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => Delay17No9_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg246_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay19No6_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg262_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg293_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg34_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg56_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg48_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => Delay80No3_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => Delay81No_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg254_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg265_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg259_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg268_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg258_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg218_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay63No_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay64No_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg240_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_impl_0_out,
                 Y => Delay1No42_out);

SharedReg249_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_1_cast <= SharedReg249_out;
SharedReg65_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_2_cast <= SharedReg65_out;
SharedReg187_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_3_cast <= SharedReg187_out;
SharedReg48_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_4_cast <= SharedReg48_out;
SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_5_cast <= SharedReg32_out;
SharedReg34_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_6_cast <= SharedReg34_out;
Delay34No1_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_7_cast <= Delay34No1_out;
SharedReg41_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_8_cast <= SharedReg41_out;
SharedReg70_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_9_cast <= SharedReg70_out;
SharedReg203_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_10_cast <= SharedReg203_out;
SharedReg203_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_11_cast <= SharedReg203_out;
SharedReg208_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_12_cast <= SharedReg208_out;
SharedReg187_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_13_cast <= SharedReg187_out;
SharedReg59_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_14_cast <= SharedReg59_out;
SharedReg33_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_15_cast <= SharedReg33_out;
SharedReg167_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_16_cast <= SharedReg167_out;
Delay44No1_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_17_cast <= Delay44No1_out;
SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_18_cast <= SharedReg32_out;
SharedReg205_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_19_cast <= SharedReg205_out;
SharedReg39_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_20_cast <= SharedReg39_out;
SharedReg49_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_21_cast <= SharedReg49_out;
SharedReg291_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_22_cast <= SharedReg291_out;
SharedReg299_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_23_cast <= SharedReg299_out;
SharedReg285_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_24_cast <= SharedReg285_out;
SharedReg52_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_25_cast <= SharedReg52_out;
SharedReg54_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_26_cast <= SharedReg54_out;
SharedReg48_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_27_cast <= SharedReg48_out;
SharedReg165_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_28_cast <= SharedReg165_out;
   MUX_Product21_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg249_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg65_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg203_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg208_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg187_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg59_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg33_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg167_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => Delay44No1_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg205_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg39_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg187_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg49_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg291_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg299_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg285_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg52_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg54_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg48_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg165_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg48_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg34_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay34No1_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg41_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg70_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg203_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Subtract2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_impl_out,
                 X => Delay1No44_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast);

SharedReg154_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg154_out;
SharedReg130_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
SharedReg151_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg151_out;
SharedReg141_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg141_out;
SharedReg_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg_out;
SharedReg176_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg176_out;
SharedReg97_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg97_out;
SharedReg3_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg3_out;
SharedReg158_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg158_out;
SharedReg113_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg113_out;
SharedReg100_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg100_out;
SharedReg129_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg129_out;
SharedReg181_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg181_out;
SharedReg110_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg110_out;
SharedReg103_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg103_out;
SharedReg109_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg109_out;
SharedReg105_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg105_out;
SharedReg96_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg96_out;
SharedReg107_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg107_out;
SharedReg154_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg154_out;
SharedReg107_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg107_out;
SharedReg176_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg176_out;
SharedReg85_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg85_out;
SharedReg150_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg150_out;
SharedReg176_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg176_out;
SharedReg97_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg97_out;
SharedReg155_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg155_out;
SharedReg96_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg96_out;
   MUX_Subtract2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg154_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg100_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg129_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg181_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg110_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg103_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg109_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg105_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg96_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg107_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg154_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg151_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg107_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg176_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg85_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg150_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg176_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg97_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg155_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg96_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg141_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg176_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg97_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg3_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg158_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg113_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_impl_0_out,
                 Y => Delay1No44_out);

SharedReg111_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg141_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg141_out;
SharedReg164_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg164_out;
SharedReg161_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg161_out;
SharedReg16_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg16_out;
SharedReg155_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg155_out;
SharedReg110_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg110_out;
SharedReg19_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg19_out;
SharedReg140_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg140_out;
SharedReg139_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg139_out;
SharedReg133_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg133_out;
SharedReg126_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg126_out;
SharedReg223_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg223_out;
Delay33No1_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_14_cast <= Delay33No1_out;
SharedReg136_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg136_out;
SharedReg130_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg130_out;
SharedReg112_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg112_out;
SharedReg104_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg104_out;
SharedReg101_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg101_out;
SharedReg176_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg176_out;
SharedReg108_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg108_out;
SharedReg96_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg96_out;
SharedReg33_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg33_out;
SharedReg130_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg130_out;
SharedReg221_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg221_out;
SharedReg141_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg141_out;
SharedReg108_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg108_out;
SharedReg108_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg108_out;
   MUX_Subtract2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg141_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg133_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg126_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg223_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay33No1_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg136_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg130_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg112_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg104_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg101_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg176_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg164_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg108_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg96_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg33_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg130_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg221_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg141_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg108_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg108_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg161_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg16_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg155_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg110_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg19_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg140_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg139_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Product13_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Product13_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Product13_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product13_impl_out,
                 X => Delay1No46_out_to_Product13_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Product13_impl_parent_implementedSystem_port_1_cast);

SharedReg79_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast <= SharedReg79_out;
SharedReg82_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast <= SharedReg82_out;
SharedReg262_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_3_cast <= SharedReg262_out;
SharedReg32_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_4_cast <= SharedReg32_out;
SharedReg268_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_5_cast <= SharedReg268_out;
SharedReg266_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_6_cast <= SharedReg266_out;
Delay62No_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_7_cast <= Delay62No_out;
SharedReg209_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_8_cast <= SharedReg209_out;
SharedReg52_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_9_cast <= SharedReg52_out;
SharedReg241_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_10_cast <= SharedReg241_out;
SharedReg277_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_11_cast <= SharedReg277_out;
SharedReg208_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_12_cast <= SharedReg208_out;
Delay96No_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_13_cast <= Delay96No_out;
Delay69No2_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_14_cast <= Delay69No2_out;
Delay14No5_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_15_cast <= Delay14No5_out;
SharedReg207_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_16_cast <= SharedReg207_out;
SharedReg302_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_17_cast <= SharedReg302_out;
Delay17No10_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_18_cast <= Delay17No10_out;
SharedReg247_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_19_cast <= SharedReg247_out;
SharedReg39_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_20_cast <= SharedReg39_out;
SharedReg189_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_21_cast <= SharedReg189_out;
Delay105No_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_22_cast <= Delay105No_out;
Delay78No3_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_23_cast <= Delay78No3_out;
SharedReg290_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_24_cast <= SharedReg290_out;
Delay80No_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_25_cast <= Delay80No_out;
Delay81No1_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_26_cast <= Delay81No1_out;
SharedReg254_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_27_cast <= SharedReg254_out;
SharedReg219_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_28_cast <= SharedReg219_out;
   MUX_Product13_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg79_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg82_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg277_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg208_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay96No_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay69No2_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay14No5_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg207_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg302_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => Delay17No10_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg247_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg39_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg262_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg189_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay105No_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => Delay78No3_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg290_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => Delay80No_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => Delay81No1_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg254_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg219_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg32_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg268_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg266_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay62No_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg209_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg52_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg241_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product13_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_impl_0_out,
                 Y => Delay1No46_out);

SharedReg261_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast <= SharedReg261_out;
SharedReg251_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast <= SharedReg251_out;
SharedReg119_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_3_cast <= SharedReg119_out;
SharedReg259_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_4_cast <= SharedReg259_out;
SharedReg35_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_5_cast <= SharedReg35_out;
SharedReg32_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_6_cast <= SharedReg32_out;
SharedReg40_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_7_cast <= SharedReg40_out;
Delay63No1_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_8_cast <= Delay63No1_out;
SharedReg255_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_9_cast <= SharedReg255_out;
SharedReg203_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_10_cast <= SharedReg203_out;
SharedReg203_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_11_cast <= SharedReg203_out;
Delay11No20_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_12_cast <= Delay11No20_out;
SharedReg77_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_13_cast <= SharedReg77_out;
SharedReg48_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_14_cast <= SharedReg48_out;
SharedReg32_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_15_cast <= SharedReg32_out;
Delay15No2_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_16_cast <= Delay15No2_out;
SharedReg117_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_17_cast <= SharedReg117_out;
SharedReg187_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_18_cast <= SharedReg187_out;
SharedReg204_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_19_cast <= SharedReg204_out;
Delay19No7_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_20_cast <= Delay19No7_out;
SharedReg295_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_21_cast <= SharedReg295_out;
SharedReg35_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_22_cast <= SharedReg35_out;
SharedReg68_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_23_cast <= SharedReg68_out;
SharedReg36_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_24_cast <= SharedReg36_out;
SharedReg49_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_25_cast <= SharedReg49_out;
SharedReg32_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_26_cast <= SharedReg32_out;
SharedReg62_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_27_cast <= SharedReg62_out;
SharedReg265_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_28_cast <= SharedReg265_out;
   MUX_Product13_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg261_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg251_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg203_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay11No20_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg77_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg48_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg32_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay15No2_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg117_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg187_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg204_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay19No7_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg119_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg295_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg35_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg68_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg36_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg49_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg32_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg62_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg265_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg259_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg35_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg32_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg40_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay63No1_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg255_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg203_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product13_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Product23_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Product23_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Product23_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_impl_out,
                 X => Delay1No48_out_to_Product23_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Product23_impl_parent_implementedSystem_port_1_cast);

SharedReg270_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_1_cast <= SharedReg270_out;
SharedReg252_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_2_cast <= SharedReg252_out;
SharedReg263_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_3_cast <= SharedReg263_out;
Delay59No1_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_4_cast <= Delay59No1_out;
SharedReg269_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_5_cast <= SharedReg269_out;
SharedReg282_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_6_cast <= SharedReg282_out;
SharedReg279_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_7_cast <= SharedReg279_out;
Delay35No2_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_8_cast <= Delay35No2_out;
SharedReg256_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_9_cast <= SharedReg256_out;
SharedReg324_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_10_cast <= SharedReg324_out;
SharedReg300_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_11_cast <= SharedReg300_out;
Delay39No_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_12_cast <= Delay39No_out;
Delay96No2_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_13_cast <= Delay96No2_out;
SharedReg316_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_14_cast <= SharedReg316_out;
Delay14No6_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_15_cast <= Delay14No6_out;
Delay43No1_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_16_cast <= Delay43No1_out;
SharedReg302_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_17_cast <= SharedReg302_out;
SharedReg237_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_18_cast <= SharedReg237_out;
SharedReg278_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_19_cast <= SharedReg278_out;
Delay103No2_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_20_cast <= Delay103No2_out;
SharedReg298_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_21_cast <= SharedReg298_out;
SharedReg35_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_22_cast <= SharedReg35_out;
SharedReg67_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_23_cast <= SharedReg67_out;
Delay79No6_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_24_cast <= Delay79No6_out;
Delay80No1_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_25_cast <= Delay80No1_out;
SharedReg73_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_26_cast <= SharedReg73_out;
Delay54No3_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_27_cast <= Delay54No3_out;
Delay55No6_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_28_cast <= Delay55No6_out;
   MUX_Product23_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg270_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg252_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg300_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay39No_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay96No2_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg316_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay14No6_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay43No1_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg302_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg237_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg278_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay103No2_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg263_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg298_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg35_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg67_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => Delay79No6_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => Delay80No1_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg73_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => Delay54No3_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => Delay55No6_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => Delay59No1_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg269_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg282_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg279_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay35No2_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg256_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg324_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product23_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_impl_0_out,
                 Y => Delay1No48_out);

SharedReg203_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_1_cast <= SharedReg203_out;
SharedReg35_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_2_cast <= SharedReg35_out;
SharedReg187_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_3_cast <= SharedReg187_out;
SharedReg65_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_4_cast <= SharedReg65_out;
SharedReg32_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_5_cast <= SharedReg32_out;
SharedReg203_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_6_cast <= SharedReg203_out;
SharedReg75_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_7_cast <= SharedReg75_out;
SharedReg189_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_8_cast <= SharedReg189_out;
SharedReg34_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_9_cast <= SharedReg34_out;
SharedReg117_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_10_cast <= SharedReg117_out;
SharedReg48_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_11_cast <= SharedReg48_out;
SharedReg38_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_12_cast <= SharedReg38_out;
SharedReg218_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_13_cast <= SharedReg218_out;
SharedReg187_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_14_cast <= SharedReg187_out;
SharedReg86_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_15_cast <= SharedReg86_out;
Delay28No2_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_16_cast <= Delay28No2_out;
SharedReg165_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_17_cast <= SharedReg165_out;
SharedReg169_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_18_cast <= SharedReg169_out;
SharedReg65_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_19_cast <= SharedReg65_out;
SharedReg196_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_20_cast <= SharedReg196_out;
SharedReg55_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_21_cast <= SharedReg55_out;
Delay105No1_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_22_cast <= Delay105No1_out;
SharedReg305_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_23_cast <= SharedReg305_out;
SharedReg65_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_24_cast <= SharedReg65_out;
SharedReg33_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_25_cast <= SharedReg33_out;
SharedReg313_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_26_cast <= SharedReg313_out;
SharedReg48_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_27_cast <= SharedReg48_out;
SharedReg201_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_28_cast <= SharedReg201_out;
   MUX_Product23_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg203_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg35_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg48_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg38_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg218_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg187_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg86_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay28No2_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg165_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg169_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg65_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg196_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg187_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg55_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay105No1_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg305_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg65_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg33_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg313_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg48_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg201_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg65_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg32_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg203_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg75_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg189_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg34_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg117_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product23_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Product33_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Product33_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Product33_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_impl_out,
                 X => Delay1No50_out_to_Product33_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Product33_impl_parent_implementedSystem_port_1_cast);

SharedReg203_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_1_cast <= SharedReg203_out;
SharedReg35_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_2_cast <= SharedReg35_out;
SharedReg119_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_3_cast <= SharedReg119_out;
Delay59No2_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_4_cast <= Delay59No2_out;
SharedReg35_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_5_cast <= SharedReg35_out;
SharedReg283_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_6_cast <= SharedReg283_out;
SharedReg61_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_7_cast <= SharedReg61_out;
SharedReg207_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_8_cast <= SharedReg207_out;
Delay64No1_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_9_cast <= Delay64No1_out;
SharedReg324_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_10_cast <= SharedReg324_out;
SharedReg48_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_11_cast <= SharedReg48_out;
SharedReg257_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_12_cast <= SharedReg257_out;
Delay96No1_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_13_cast <= Delay96No1_out;
Delay69No5_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_14_cast <= Delay69No5_out;
SharedReg86_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_15_cast <= SharedReg86_out;
SharedReg296_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_16_cast <= SharedReg296_out;
SharedReg303_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_17_cast <= SharedReg303_out;
SharedReg187_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_18_cast <= SharedReg187_out;
SharedReg322_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_19_cast <= SharedReg322_out;
Delay103No3_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_20_cast <= Delay103No3_out;
SharedReg304_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_21_cast <= SharedReg304_out;
Delay77No2_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_22_cast <= Delay77No2_out;
SharedReg289_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_23_cast <= SharedReg289_out;
SharedReg288_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_24_cast <= SharedReg288_out;
Delay80No4_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_25_cast <= Delay80No4_out;
SharedReg206_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_26_cast <= SharedReg206_out;
Delay54No4_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_27_cast <= Delay54No4_out;
SharedReg274_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_28_cast <= SharedReg274_out;
   MUX_Product33_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg203_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg35_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg48_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg257_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay96No1_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay69No5_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg86_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg296_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg303_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg187_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg322_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay103No3_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg119_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg304_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay77No2_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg289_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg288_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => Delay80No4_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg206_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => Delay54No4_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg274_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => Delay59No2_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg35_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg283_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg61_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg207_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay64No1_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg324_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_impl_0_out,
                 Y => Delay1No50_out);

SharedReg271_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_1_cast <= SharedReg271_out;
SharedReg253_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_2_cast <= SharedReg253_out;
SharedReg263_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_3_cast <= SharedReg263_out;
SharedReg65_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_4_cast <= SharedReg65_out;
SharedReg269_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_5_cast <= SharedReg269_out;
SharedReg187_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_6_cast <= SharedReg187_out;
SharedReg279_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_7_cast <= SharedReg279_out;
Delay35No1_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_8_cast <= Delay35No1_out;
SharedReg209_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_9_cast <= SharedReg209_out;
SharedReg166_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_10_cast <= SharedReg166_out;
SharedReg301_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_11_cast <= SharedReg301_out;
SharedReg37_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_12_cast <= SharedReg37_out;
SharedReg217_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_13_cast <= SharedReg217_out;
SharedReg187_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_14_cast <= SharedReg187_out;
Delay14No7_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_15_cast <= Delay14No7_out;
SharedReg187_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_16_cast <= SharedReg187_out;
SharedReg117_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_17_cast <= SharedReg117_out;
SharedReg237_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_18_cast <= SharedReg237_out;
SharedReg67_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_19_cast <= SharedReg67_out;
SharedReg191_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_20_cast <= SharedReg191_out;
SharedReg65_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_21_cast <= SharedReg65_out;
SharedReg51_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_22_cast <= SharedReg51_out;
SharedReg205_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_23_cast <= SharedReg205_out;
SharedReg206_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_24_cast <= SharedReg206_out;
SharedReg66_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_25_cast <= SharedReg66_out;
SharedReg317_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_26_cast <= SharedReg317_out;
SharedReg63_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_27_cast <= SharedReg63_out;
SharedReg209_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_28_cast <= SharedReg209_out;
   MUX_Product33_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg271_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg253_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg301_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg37_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg217_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg187_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay14No7_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg187_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg117_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg237_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg67_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg191_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg263_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg65_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg51_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg205_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg206_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg66_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg317_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg63_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg209_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg65_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg269_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg187_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg279_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay35No1_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg209_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg166_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Subtract4_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Subtract4_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Subtract4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_impl_out,
                 X => Delay1No52_out_to_Subtract4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Subtract4_impl_parent_implementedSystem_port_1_cast);

SharedReg65_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg65_out;
SharedReg176_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg176_out;
SharedReg128_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg128_out;
SharedReg1_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1_out;
SharedReg117_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg117_out;
SharedReg162_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg162_out;
SharedReg123_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg123_out;
SharedReg57_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg57_out;
Delay8No1_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_9_cast <= Delay8No1_out;
SharedReg143_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg143_out;
Delay28No3_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_11_cast <= Delay28No3_out;
SharedReg95_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg95_out;
Delay12No_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_13_cast <= Delay12No_out;
SharedReg141_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg141_out;
SharedReg225_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg225_out;
SharedReg100_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg100_out;
SharedReg154_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg154_out;
SharedReg141_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg141_out;
SharedReg152_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg152_out;
SharedReg221_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg221_out;
SharedReg113_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg113_out;
SharedReg110_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg110_out;
SharedReg188_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg188_out;
SharedReg181_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg181_out;
SharedReg117_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg117_out;
SharedReg65_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg65_out;
SharedReg130_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg130_out;
SharedReg98_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg98_out;
   MUX_Subtract4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg65_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg176_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay28No3_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg95_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay12No_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg141_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg225_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg100_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg154_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg141_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg152_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg221_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg128_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg113_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg110_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg188_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg181_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg117_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg65_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg130_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg98_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg117_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg162_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg123_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg57_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay8No1_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg143_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_impl_0_out,
                 Y => Delay1No52_out);

SharedReg82_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg82_out;
SharedReg221_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg221_out;
SharedReg117_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg117_out;
SharedReg17_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg17_out;
SharedReg165_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg165_out;
SharedReg137_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg137_out;
SharedReg117_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg117_out;
SharedReg82_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg82_out;
Delay8No3_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_9_cast <= Delay8No3_out;
SharedReg133_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg133_out;
SharedReg177_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg177_out;
SharedReg92_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg92_out;
Delay12No5_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_13_cast <= Delay12No5_out;
SharedReg221_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg221_out;
SharedReg227_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg227_out;
SharedReg99_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg99_out;
SharedReg182_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg182_out;
SharedReg160_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg160_out;
SharedReg159_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg159_out;
SharedReg138_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg138_out;
SharedReg131_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg131_out;
SharedReg154_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg154_out;
SharedReg118_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg118_out;
SharedReg157_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg157_out;
SharedReg165_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg165_out;
SharedReg82_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg82_out;
SharedReg141_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg141_out;
SharedReg97_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg97_out;
   MUX_Subtract4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg82_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg221_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg177_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg92_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay12No5_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg221_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg227_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg99_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg182_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg160_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg159_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg138_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg117_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg131_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg154_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg118_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg157_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg165_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg82_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg141_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg97_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg17_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg165_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg137_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg117_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg82_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay8No3_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg133_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Product7_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Product7_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Product7_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product7_impl_out,
                 X => Delay1No54_out_to_Product7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Product7_impl_parent_implementedSystem_port_1_cast);

SharedReg220_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg220_out;
SharedReg165_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg165_out;
SharedReg195_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg195_out;
SharedReg189_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg189_out;
SharedReg275_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg275_out;
SharedReg238_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg238_out;
SharedReg244_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg244_out;
Delay60No_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_8_cast <= Delay60No_out;
SharedReg260_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg260_out;
Delay57No3_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_10_cast <= Delay57No3_out;
SharedReg272_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg272_out;
SharedReg281_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg281_out;
SharedReg288_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg288_out;
Delay103No_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_14_cast <= Delay103No_out;
Delay34No4_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_15_cast <= Delay34No4_out;
SharedReg307_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg307_out;
SharedReg308_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg308_out;
Delay78No6_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_18_cast <= Delay78No6_out;
Delay81No3_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_19_cast <= Delay81No3_out;
SharedReg314_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg314_out;
SharedReg318_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg318_out;
SharedReg320_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg320_out;
Delay42No_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_23_cast <= Delay42No_out;
SharedReg325_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg325_out;
Delay18No10_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_25_cast <= Delay18No10_out;
SharedReg326_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg326_out;
   MUX_Product7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_26_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg220_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg165_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg272_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg281_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg288_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay103No_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay34No4_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg307_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg308_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => Delay78No6_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => Delay81No3_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg314_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg195_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg318_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg320_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => Delay42No_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg325_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => Delay18No10_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg326_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_3 => SharedReg189_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg275_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg238_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg244_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay60No_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg260_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay57No3_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product7_impl_0_LUT_out,
                 oMux => MUX_Product7_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product7_impl_0_out,
                 Y => Delay1No54_out);

SharedReg78_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg78_out;
SharedReg43_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg43_out;
SharedReg65_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg65_out;
SharedReg32_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg32_out;
SharedReg64_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg64_out;
SharedReg117_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg117_out;
SharedReg166_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg166_out;
SharedReg117_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg117_out;
SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg187_out;
SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg187_out;
SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg187_out;
SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg187_out;
SharedReg203_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg203_out;
Delay30No2_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_14_cast <= Delay30No2_out;
SharedReg205_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg205_out;
SharedReg190_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg190_out;
SharedReg205_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg205_out;
SharedReg204_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg204_out;
SharedReg203_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg203_out;
SharedReg212_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg212_out;
SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg187_out;
SharedReg204_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg204_out;
Delay61No_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_23_cast <= Delay61No_out;
SharedReg297_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg297_out;
SharedReg303_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg303_out;
Delay80No5_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_26_cast <= Delay80No5_out;
   MUX_Product7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_26_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg78_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg43_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg203_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay30No2_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg205_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg190_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg205_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg204_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg203_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg212_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg65_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg204_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => Delay61No_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg297_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg303_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => Delay80No5_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_3 => SharedReg32_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg64_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg117_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg166_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg117_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg187_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product7_impl_1_LUT_out,
                 oMux => MUX_Product7_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product7_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Subtract17_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Subtract17_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Subtract17_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract17_impl_out,
                 X => Delay1No56_out_to_Subtract17_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Subtract17_impl_parent_implementedSystem_port_1_cast);

SharedReg117_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg58_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_2_cast <= SharedReg58_out;
SharedReg94_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_3_cast <= SharedReg94_out;
SharedReg117_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_4_cast <= SharedReg117_out;
SharedReg193_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_5_cast <= SharedReg193_out;
SharedReg65_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_6_cast <= SharedReg65_out;
SharedReg173_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_7_cast <= SharedReg173_out;
SharedReg10_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_8_cast <= SharedReg10_out;
SharedReg200_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_9_cast <= SharedReg200_out;
SharedReg111_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_10_cast <= SharedReg111_out;
SharedReg129_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_11_cast <= SharedReg129_out;
SharedReg7_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_12_cast <= SharedReg7_out;
Delay12No2_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_13_cast <= Delay12No2_out;
SharedReg83_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_14_cast <= SharedReg83_out;
SharedReg54_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_15_cast <= SharedReg54_out;
SharedReg231_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_16_cast <= SharedReg231_out;
SharedReg185_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_17_cast <= SharedReg185_out;
SharedReg50_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_18_cast <= SharedReg50_out;
SharedReg176_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_19_cast <= SharedReg176_out;
SharedReg131_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_20_cast <= SharedReg131_out;
SharedReg130_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_21_cast <= SharedReg130_out;
SharedReg91_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_22_cast <= SharedReg91_out;
SharedReg127_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_23_cast <= SharedReg127_out;
SharedReg165_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_24_cast <= SharedReg165_out;
SharedReg118_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_25_cast <= SharedReg118_out;
SharedReg171_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_26_cast <= SharedReg171_out;
SharedReg165_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_27_cast <= SharedReg165_out;
SharedReg51_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_28_cast <= SharedReg51_out;
   MUX_Subtract17_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg58_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg129_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg7_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay12No2_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg83_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg54_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg231_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg185_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg50_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg176_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg131_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg94_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg130_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg91_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg127_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg165_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg118_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg171_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg165_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg51_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg117_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg193_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg65_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg173_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg10_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg200_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg111_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract17_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract17_impl_0_out,
                 Y => Delay1No56_out);

SharedReg165_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_1_cast <= SharedReg165_out;
Delay44No_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_2_cast <= Delay44No_out;
SharedReg82_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_3_cast <= SharedReg82_out;
SharedReg165_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_4_cast <= SharedReg165_out;
SharedReg210_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_5_cast <= SharedReg210_out;
SharedReg82_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_6_cast <= SharedReg82_out;
SharedReg165_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_7_cast <= SharedReg165_out;
SharedReg26_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_8_cast <= SharedReg26_out;
SharedReg117_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_9_cast <= SharedReg117_out;
SharedReg156_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_10_cast <= SharedReg156_out;
Delay24No3_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_11_cast <= Delay24No3_out;
SharedReg23_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_12_cast <= SharedReg23_out;
Delay12No7_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_13_cast <= Delay12No7_out;
SharedReg82_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_14_cast <= SharedReg82_out;
SharedReg71_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_15_cast <= SharedReg71_out;
SharedReg222_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_16_cast <= SharedReg222_out;
Delay29No17_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_17_cast <= Delay29No17_out;
SharedReg67_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_18_cast <= SharedReg67_out;
SharedReg221_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_19_cast <= SharedReg221_out;
SharedReg157_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_20_cast <= SharedReg157_out;
SharedReg176_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_21_cast <= SharedReg176_out;
SharedReg65_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_22_cast <= SharedReg65_out;
SharedReg167_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_23_cast <= SharedReg167_out;
SharedReg187_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_24_cast <= SharedReg187_out;
SharedReg202_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_25_cast <= SharedReg202_out;
SharedReg165_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_26_cast <= SharedReg165_out;
SharedReg120_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_27_cast <= SharedReg120_out;
SharedReg85_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_28_cast <= SharedReg85_out;
   MUX_Subtract17_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg165_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay44No_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay24No3_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg23_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay12No7_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg82_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg71_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg222_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => Delay29No17_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg67_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg221_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg157_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg82_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg176_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg65_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg167_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg187_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg202_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg165_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg120_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg85_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg165_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg210_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg82_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg165_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg26_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg117_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg156_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract17_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract17_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Subtract20_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Subtract20_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Subtract20_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract20_impl_out,
                 X => Delay1No58_out_to_Subtract20_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Subtract20_impl_parent_implementedSystem_port_1_cast);

SharedReg48_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_1_cast <= SharedReg48_out;
SharedReg13_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg6_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_3_cast <= SharedReg6_out;
SharedReg82_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_4_cast <= SharedReg82_out;
SharedReg8_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_5_cast <= SharedReg8_out;
SharedReg12_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_6_cast <= SharedReg12_out;
Delay6No_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_7_cast <= Delay6No_out;
Delay7No3_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_8_cast <= Delay7No3_out;
SharedReg65_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_9_cast <= SharedReg65_out;
SharedReg109_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_10_cast <= SharedReg109_out;
SharedReg165_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_11_cast <= SharedReg165_out;
SharedReg15_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_12_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_13_cast <= SharedReg14_out;
SharedReg120_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_14_cast <= SharedReg120_out;
SharedReg117_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_15_cast <= SharedReg117_out;
SharedReg117_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_16_cast <= SharedReg117_out;
SharedReg60_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_17_cast <= SharedReg60_out;
SharedReg82_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_18_cast <= SharedReg82_out;
SharedReg66_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_19_cast <= SharedReg66_out;
SharedReg117_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_20_cast <= SharedReg117_out;
SharedReg162_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_21_cast <= SharedReg162_out;
SharedReg125_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_22_cast <= SharedReg125_out;
SharedReg65_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_23_cast <= SharedReg65_out;
SharedReg82_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_24_cast <= SharedReg82_out;
SharedReg32_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_25_cast <= SharedReg32_out;
SharedReg117_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_26_cast <= SharedReg117_out;
SharedReg65_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_27_cast <= SharedReg65_out;
SharedReg82_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_28_cast <= SharedReg82_out;
   MUX_Subtract20_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg48_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg165_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg15_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg14_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg120_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg117_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg117_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg60_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg82_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg66_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg117_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg6_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg162_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg125_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg65_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg82_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg32_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg117_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg65_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg82_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg82_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg8_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg12_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay6No_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay7No3_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg65_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg109_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract20_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_impl_0_out,
                 Y => Delay1No58_out);

SharedReg69_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_1_cast <= SharedReg69_out;
SharedReg29_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_2_cast <= SharedReg29_out;
SharedReg22_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_3_cast <= SharedReg22_out;
SharedReg90_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_4_cast <= SharedReg90_out;
SharedReg24_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_5_cast <= SharedReg24_out;
SharedReg28_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_6_cast <= SharedReg28_out;
Delay6No2_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_7_cast <= Delay6No2_out;
Delay7No7_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_8_cast <= Delay7No7_out;
SharedReg82_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_9_cast <= SharedReg82_out;
SharedReg155_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_10_cast <= SharedReg155_out;
SharedReg126_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_11_cast <= SharedReg126_out;
SharedReg31_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_12_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_13_cast <= SharedReg30_out;
SharedReg117_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_14_cast <= SharedReg117_out;
SharedReg165_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_15_cast <= SharedReg165_out;
SharedReg204_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_16_cast <= SharedReg204_out;
SharedReg76_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_17_cast <= SharedReg76_out;
SharedReg85_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_18_cast <= SharedReg85_out;
SharedReg84_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_19_cast <= SharedReg84_out;
SharedReg165_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_20_cast <= SharedReg165_out;
SharedReg230_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_21_cast <= SharedReg230_out;
SharedReg165_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_22_cast <= SharedReg165_out;
SharedReg82_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_23_cast <= SharedReg82_out;
SharedReg89_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_24_cast <= SharedReg89_out;
SharedReg94_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_25_cast <= SharedReg94_out;
SharedReg192_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_26_cast <= SharedReg192_out;
SharedReg87_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_27_cast <= SharedReg87_out;
SharedReg53_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_28_cast <= SharedReg53_out;
   MUX_Subtract20_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg126_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg31_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg30_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg117_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg165_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg204_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg76_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg85_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg84_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg165_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg22_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg230_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg165_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg82_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg89_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg94_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg192_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg87_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg53_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg90_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg24_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg28_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay6No2_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay7No7_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg82_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg155_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract20_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Product220_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Product220_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Product220_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product220_impl_out,
                 X => Delay1No60_out_to_Product220_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Product220_impl_parent_implementedSystem_port_1_cast);

SharedReg81_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_1_cast <= SharedReg81_out;
SharedReg80_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_2_cast <= SharedReg80_out;
SharedReg166_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_3_cast <= SharedReg166_out;
SharedReg117_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_4_cast <= SharedReg117_out;
SharedReg187_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_5_cast <= SharedReg187_out;
SharedReg209_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_6_cast <= SharedReg209_out;
SharedReg203_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_7_cast <= SharedReg203_out;
SharedReg188_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_8_cast <= SharedReg188_out;
SharedReg213_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_9_cast <= SharedReg213_out;
SharedReg245_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_10_cast <= SharedReg245_out;
Delay57No4_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_11_cast <= Delay57No4_out;
SharedReg273_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_12_cast <= SharedReg273_out;
Delay59No3_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_13_cast <= Delay59No3_out;
SharedReg280_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_14_cast <= SharedReg280_out;
SharedReg294_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_15_cast <= SharedReg294_out;
Delay103No1_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_16_cast <= Delay103No1_out;
SharedReg306_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_17_cast <= SharedReg306_out;
SharedReg312_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_18_cast <= SharedReg312_out;
Delay82No_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_19_cast <= Delay82No_out;
Delay97No_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_20_cast <= Delay97No_out;
Delay80No6_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_21_cast <= Delay80No6_out;
Delay16No8_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_22_cast <= Delay16No8_out;
SharedReg319_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_23_cast <= SharedReg319_out;
SharedReg321_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_24_cast <= SharedReg321_out;
SharedReg323_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_25_cast <= SharedReg323_out;
Delay18No11_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_26_cast <= Delay18No11_out;
   MUX_Product220_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_26_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg81_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg80_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay57No4_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg273_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay59No3_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg280_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg294_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay103No1_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg306_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg312_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => Delay82No_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay97No_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg166_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => Delay80No6_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay16No8_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg319_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg321_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg323_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => Delay18No11_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_26_cast,
                 iS_3 => SharedReg117_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg187_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg209_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg203_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg188_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg213_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg245_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product220_impl_0_LUT_out,
                 oMux => MUX_Product220_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product220_impl_0_out,
                 Y => Delay1No60_out);

SharedReg33_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_1_cast <= SharedReg33_out;
SharedReg72_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_2_cast <= SharedReg72_out;
SharedReg33_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_3_cast <= SharedReg33_out;
SharedReg34_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_4_cast <= SharedReg34_out;
SharedReg32_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_5_cast <= SharedReg32_out;
SharedReg60_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_6_cast <= SharedReg60_out;
SharedReg166_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_7_cast <= SharedReg166_out;
SharedReg187_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_8_cast <= SharedReg187_out;
SharedReg205_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_9_cast <= SharedReg205_out;
SharedReg191_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_10_cast <= SharedReg191_out;
SharedReg203_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_11_cast <= SharedReg203_out;
SharedReg207_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_12_cast <= SharedReg207_out;
SharedReg187_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_13_cast <= SharedReg187_out;
Delay31No_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_14_cast <= Delay31No_out;
SharedReg214_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_15_cast <= SharedReg214_out;
SharedReg275_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_16_cast <= SharedReg275_out;
SharedReg187_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_17_cast <= SharedReg187_out;
SharedReg203_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_18_cast <= SharedReg203_out;
Delay60No1_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_19_cast <= Delay60No1_out;
Delay79No4_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_20_cast <= Delay79No4_out;
SharedReg309_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_21_cast <= SharedReg309_out;
SharedReg315_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_22_cast <= SharedReg315_out;
Delay38No_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_23_cast <= Delay38No_out;
Delay42No1_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_24_cast <= Delay42No1_out;
SharedReg325_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_25_cast <= SharedReg325_out;
SharedReg327_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_26_cast <= SharedReg327_out;
   MUX_Product220_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_26_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg33_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg203_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg207_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg187_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay31No_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg214_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg275_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg187_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg203_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => Delay60No1_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay79No4_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg33_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg309_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg315_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => Delay38No_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => Delay42No1_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg325_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg327_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_26_cast,
                 iS_3 => SharedReg34_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg32_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg60_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg166_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg187_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg205_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg191_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product220_impl_1_LUT_out,
                 oMux => MUX_Product220_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product220_impl_1_out,
                 Y => Delay1No61_out);
   Constant2_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant2_impl_out);
   Constant11_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant11_impl_out);
   Constant3_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant3_impl_out);
   Constant12_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant12_impl_out);
   Constant4_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant4_impl_out);
   Constant13_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant13_impl_out);
   Constant5_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant5_impl_out);
   Constant14_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant14_impl_out);
   Constant6_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant6_impl_out);
   Constant15_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant15_impl_out);
   Constant7_impl_instance: Constant_float_8_23_cosn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant7_impl_out);
   Constant16_impl_instance: Constant_float_8_23_sinn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant16_impl_out);
   Constant8_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant8_impl_out);
   Constant17_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant17_impl_out);
   Constant9_impl_instance: Constant_float_8_23_cosn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant9_impl_out);
   Constant18_impl_instance: Constant_float_8_23_sinn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant18_impl_out);
   Constant10_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant10_impl_out);
   Constant19_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant19_impl_out);
   Constant20_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant20_impl_out);
   Constant110_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant110_impl_out);
   Constant21_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant21_impl_out);
   Constant111_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant111_impl_out);
   Constant22_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant22_impl_out);
   Constant112_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant112_impl_out);
   Constant23_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant23_impl_out);
   Constant113_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant113_impl_out);
   Constant24_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant24_impl_out);
   Constant114_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant114_impl_out);
   Constant25_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant25_impl_out);
   Constant115_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant115_impl_out);
   Constant26_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant26_impl_out);
   Constant116_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant116_impl_out);
   Constant27_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant27_impl_out);
   Constant117_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant117_impl_out);
   Constant28_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant28_impl_out);
   Constant118_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant118_impl_out);
   Constant29_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant29_impl_out);
   Constant119_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant119_impl_out);
   Constant30_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant30_impl_out);
   Constant120_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant120_impl_out);
   Constant31_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant31_impl_out);
   Constant121_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant121_impl_out);
   Constant32_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant32_impl_out);
   Constant122_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant122_impl_out);
   Constant33_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant33_impl_out);
   Constant123_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant123_impl_out);
   Constant34_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant34_impl_out);
   Constant124_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant124_impl_out);
   Constant35_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant35_impl_out);
   Constant125_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant125_impl_out);
   Constant36_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant36_impl_out);
   Constant126_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant126_impl_out);
   Constant37_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant37_impl_out);
   Constant127_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant127_impl_out);
   Constant38_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant38_impl_out);
   Constant128_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant128_impl_out);
   Constant39_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant39_impl_out);
   Constant129_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant129_impl_out);
   Constant40_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant40_impl_out);
   Constant130_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant130_impl_out);
   Constant41_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant41_impl_out);
   Constant131_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant131_impl_out);
   Constant42_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant42_impl_out);
   Constant132_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant132_impl_out);
   Constant43_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant43_impl_out);
   Constant133_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant133_impl_out);
   Constant44_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant44_impl_out);
   Constant134_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant134_impl_out);
   Constant45_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant45_impl_out);
   Constant135_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant135_impl_out);
   Constant46_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant46_impl_out);
   Constant136_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant136_impl_out);
   Constant47_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant47_impl_out);
   Constant137_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant137_impl_out);
   Constant48_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant48_impl_out);
   Constant138_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant138_impl_out);
   Constant49_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant49_impl_out);
   Constant139_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant139_impl_out);
   Constant50_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant50_impl_out);
   Constant140_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant140_impl_out);
   Constant51_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant51_impl_out);
   Constant141_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant141_impl_out);
   Constant52_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant52_impl_out);
   Constant142_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant142_impl_out);
   Constant53_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant53_impl_out);
   Constant143_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant143_impl_out);
   Constant54_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant54_impl_out);
   Constant144_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant144_impl_out);
   Constant55_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant55_impl_out);
   Constant145_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant145_impl_out);
   Constant56_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant56_impl_out);
   Constant146_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant146_impl_out);
   Constant57_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant57_impl_out);
   Constant147_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant147_impl_out);
   Constant_impl_instance: Constant_float_8_23_cosnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_impl_out);
   Constant1_impl_instance: Constant_float_8_23_sinnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_impl_out);

   Delay8No_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg_out,
                 Y => Delay8No_out);

   Delay7No_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1_out,
                 Y => Delay7No_out);

   Delay12No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg2_out,
                 Y => Delay12No_out);

   Delay12No1_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg3_out,
                 Y => Delay12No1_out);

   Delay8No1_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg4_out,
                 Y => Delay8No1_out);

   Delay12No2_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => Delay12No2_out);

   Delay13No_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg6_out,
                 Y => Delay13No_out);

   Delay9No_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg8_out,
                 Y => Delay9No_out);

   Delay6No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg9_out,
                 Y => Delay6No_out);

   Delay10No_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg10_out,
                 Y => Delay10No_out);

   Delay7No3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg11_out,
                 Y => Delay7No3_out);

   Delay6No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg12_out,
                 Y => Delay6No1_out);

   Delay5No3_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg13_out,
                 Y => Delay5No3_out);

   Delay8No2_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg16_out,
                 Y => Delay8No2_out);

   Delay7No4_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg17_out,
                 Y => Delay7No4_out);

   Delay12No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg18_out,
                 Y => Delay12No5_out);

   Delay12No6_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg19_out,
                 Y => Delay12No6_out);

   Delay8No3_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg20_out,
                 Y => Delay8No3_out);

   Delay12No7_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg21_out,
                 Y => Delay12No7_out);

   Delay13No1_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg22_out,
                 Y => Delay13No1_out);

   Delay9No1_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg24_out,
                 Y => Delay9No1_out);

   Delay6No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg25_out,
                 Y => Delay6No2_out);

   Delay10No1_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg26_out,
                 Y => Delay10No1_out);

   Delay7No7_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg27_out,
                 Y => Delay7No7_out);

   Delay6No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg28_out,
                 Y => Delay6No3_out);

   Delay5No7_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg29_out,
                 Y => Delay5No7_out);

   Delay28No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => Delay28No2_out);

   Delay29No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => Delay29No2_out);

   Delay33No_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => Delay33No_out);

   Delay33No1_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => Delay33No1_out);

   Delay30No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => Delay30No1_out);

   Delay44No_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => Delay44No_out);

   Delay28No3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => Delay28No3_out);

   Delay24No3_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => Delay24No3_out);

   Delay29No15_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => Delay29No15_out);

   Delay29No17_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => Delay29No17_out);

   Delay30No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => Delay30No2_out);

   Delay31No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => Delay31No_out);

   Delay34No_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => Delay34No_out);

   Delay37No_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => Delay37No_out);

   Delay17No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => Delay17No9_out);

   Delay44No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => Delay44No1_out);

   Delay17No10_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => Delay17No10_out);

   Delay18No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => Delay18No5_out);

   Delay17No14_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => Delay17No14_out);

   Delay11No17_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => Delay11No17_out);

   Delay15No2_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => Delay15No2_out);

   Delay19No5_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => Delay19No5_out);

   Delay34No1_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => Delay34No1_out);

   Delay60No_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => Delay60No_out);

   Delay60No1_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => Delay60No1_out);

   Delay35No_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => Delay35No_out);

   Delay36No_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => Delay36No_out);

   Delay57No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => Delay57No_out);

   Delay57No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => Delay57No1_out);

   Delay59No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => Delay59No_out);

   Delay64No_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => Delay64No_out);

   Delay39No_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => Delay39No_out);

   Delay54No_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => Delay54No_out);

   Delay54No3_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => Delay54No3_out);

   Delay19No6_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => Delay19No6_out);

   Delay19No7_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => Delay19No7_out);

   Delay54No4_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => Delay54No4_out);

   Delay59No1_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => Delay59No1_out);

   Delay59No2_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => Delay59No2_out);

   Delay55No_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => Delay55No_out);

   Delay63No_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => Delay63No_out);

   Delay62No_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => Delay62No_out);

   Delay57No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => Delay57No3_out);

   Delay57No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => Delay57No4_out);

   Delay64No1_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => Delay64No1_out);

   Delay63No1_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => Delay63No1_out);

   Delay59No3_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => Delay59No3_out);

   Delay11No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => Delay11No19_out);

   Delay11No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => Delay11No20_out);

   Delay43No1_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => Delay43No1_out);

   Delay55No6_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => Delay55No6_out);

   Delay35No1_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => Delay35No1_out);

   Delay35No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => Delay35No2_out);

   Delay61No_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => Delay61No_out);

   Delay80No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => Delay80No_out);

   Delay80No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => Delay80No1_out);

   Delay80No2_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => Delay80No2_out);

   Delay80No3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => Delay80No3_out);

   Delay79No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => Delay79No4_out);

   Delay80No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => Delay80No4_out);

   Delay79No6_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => Delay79No6_out);

   Delay105No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => Delay105No_out);

   Delay105No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => Delay105No1_out);

   Delay103No_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => Delay103No_out);

   Delay103No1_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => Delay103No1_out);

   Delay103No2_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => Delay103No2_out);

   Delay103No3_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => Delay103No3_out);

   Delay77No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => Delay77No2_out);

   Delay81No_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => Delay81No_out);

   Delay14No5_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => Delay14No5_out);

   Delay34No4_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => Delay34No4_out);

   Delay78No3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => Delay78No3_out);

   Delay96No_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => Delay96No_out);

   Delay96No1_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => Delay96No1_out);

   Delay80No5_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => Delay80No5_out);

   Delay78No6_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => Delay78No6_out);

   Delay96No2_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => Delay96No2_out);

   Delay69No2_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => Delay69No2_out);

   Delay81No1_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => Delay81No1_out);

   Delay82No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => Delay82No_out);

   Delay81No3_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => Delay81No3_out);

   Delay97No_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => Delay97No_out);

   Delay80No6_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => Delay80No6_out);

   Delay69No5_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => Delay69No5_out);

   Delay16No8_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => Delay16No8_out);

   Delay38No_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => Delay38No_out);

   Delay14No6_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => Delay14No6_out);

   Delay14No7_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => Delay14No7_out);

   Delay42No_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => Delay42No_out);

   Delay42No1_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => Delay42No1_out);

   Delay18No10_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => Delay18No10_out);

   Delay18No11_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => Delay18No11_out);

   MUX_Product7_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product7_impl_0_LUT_wIn_5_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_Product7_impl_0_LUT_out);

   MUX_Product7_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product7_impl_1_LUT_wIn_5_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_Product7_impl_1_LUT_out);

   MUX_Product220_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product220_impl_0_LUT_wIn_5_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_Product220_impl_0_LUT_out);

   MUX_Product220_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product220_impl_1_LUT_wIn_5_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_Product220_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_re_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_im_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_re_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_im_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_re_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_im_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_re_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_im_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_re_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_im_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_re_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_im_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_re_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_im_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_re_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_im_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_re_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_im_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_re_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_im_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_re_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_im_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_re_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_im_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_re_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_im_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_re_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_im_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_re_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_im_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_re_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_im_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_impl_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add7_impl_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_impl_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add120_impl_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_impl_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_impl_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_impl_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product13_impl_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_impl_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_impl_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_impl_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product7_impl_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract17_impl_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract20_impl_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product220_impl_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant2_impl_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant11_impl_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant3_impl_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=43 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant12_impl_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant4_impl_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant13_impl_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant5_impl_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant14_impl_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant6_impl_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant15_impl_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant7_impl_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant16_impl_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant8_impl_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant17_impl_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant9_impl_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant18_impl_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant10_impl_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant19_impl_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=58 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant20_impl_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=57 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant110_impl_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant21_impl_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant111_impl_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=54 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant22_impl_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant112_impl_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant23_impl_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant113_impl_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=33 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant24_impl_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant114_impl_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=54 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant25_impl_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant115_impl_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant26_impl_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant116_impl_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant27_impl_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=55 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant117_impl_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=33 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant28_impl_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=33 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant118_impl_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=60 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant29_impl_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=60 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant119_impl_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant30_impl_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant120_impl_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=58 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant31_impl_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=58 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant121_impl_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=55 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant32_impl_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=55 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant122_impl_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant33_impl_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant123_impl_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant34_impl_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant124_impl_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=33 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant35_impl_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant125_impl_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=33 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant36_impl_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=33 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant126_impl_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_79_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=79 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant37_impl_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_79_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=79 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant127_impl_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_77_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=77 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant38_impl_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=78 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant128_impl_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_79_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=79 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant39_impl_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=78 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant129_impl_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_79_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=79 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant40_impl_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_77_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=77 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant130_impl_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=104 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant41_impl_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=104 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant131_impl_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=99 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant42_impl_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=76 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant132_impl_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=99 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant43_impl_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=99 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant133_impl_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=76 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant44_impl_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=78 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant134_impl_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant45_impl_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant135_impl_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_100_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=100 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant46_impl_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_100_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=100 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant136_impl_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=76 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant47_impl_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=78 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant137_impl_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=78 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant48_impl_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_77_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=77 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant138_impl_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=76 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant49_impl_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=76 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant139_impl_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=69 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant50_impl_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant140_impl_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_77_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=77 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant51_impl_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=81 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant141_impl_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=69 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant52_impl_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=81 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant142_impl_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=69 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant53_impl_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant143_impl_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant54_impl_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant144_impl_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant55_impl_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant145_impl_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant56_impl_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant146_impl_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant57_impl_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant147_impl_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_impl_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_impl_out,
                 Y => SharedReg327_out);
end architecture;



library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity implementedSystem_toplevel_wrapper is
  port (
    clk, rst : in std_logic;
    shared_input : in std_logic_vector(31 downto 0);
    x0_re_enable : in std_logic;
    x0_im_enable : in std_logic;
    x1_re_enable : in std_logic;
    x1_im_enable : in std_logic;
    x2_re_enable : in std_logic;
    x2_im_enable : in std_logic;
    x3_re_enable : in std_logic;
    x3_im_enable : in std_logic;
    x4_re_enable : in std_logic;
    x4_im_enable : in std_logic;
    x5_re_enable : in std_logic;
    x5_im_enable : in std_logic;
    x6_re_enable : in std_logic;
    x6_im_enable : in std_logic;
    x7_re_enable : in std_logic;
    x7_im_enable : in std_logic;
    x8_re_enable : in std_logic;
    x8_im_enable : in std_logic;
    x9_re_enable : in std_logic;
    x9_im_enable : in std_logic;
    x10_re_enable : in std_logic;
    x10_im_enable : in std_logic;
    x11_re_enable : in std_logic;
    x11_im_enable : in std_logic;
    x12_re_enable : in std_logic;
    x12_im_enable : in std_logic;
    x13_re_enable : in std_logic;
    x13_im_enable : in std_logic;
    x14_re_enable : in std_logic;
    x14_im_enable : in std_logic;
    x15_re_enable : in std_logic;
    x15_im_enable : in std_logic;
    output_select : in std_logic_vector(4 downto 0);
    shared_output : out std_logic_vector(31 downto 0)
  );
end entity;

architecture implementedSystem_toplevel_wrapper of implementedSystem_toplevel_wrapper is
  signal x0_re_DUT_in : std_logic_vector(31 downto 0);
  signal x0_im_DUT_in : std_logic_vector(31 downto 0);
  signal x1_re_DUT_in : std_logic_vector(31 downto 0);
  signal x1_im_DUT_in : std_logic_vector(31 downto 0);
  signal x2_re_DUT_in : std_logic_vector(31 downto 0);
  signal x2_im_DUT_in : std_logic_vector(31 downto 0);
  signal x3_re_DUT_in : std_logic_vector(31 downto 0);
  signal x3_im_DUT_in : std_logic_vector(31 downto 0);
  signal x4_re_DUT_in : std_logic_vector(31 downto 0);
  signal x4_im_DUT_in : std_logic_vector(31 downto 0);
  signal x5_re_DUT_in : std_logic_vector(31 downto 0);
  signal x5_im_DUT_in : std_logic_vector(31 downto 0);
  signal x6_re_DUT_in : std_logic_vector(31 downto 0);
  signal x6_im_DUT_in : std_logic_vector(31 downto 0);
  signal x7_re_DUT_in : std_logic_vector(31 downto 0);
  signal x7_im_DUT_in : std_logic_vector(31 downto 0);
  signal x8_re_DUT_in : std_logic_vector(31 downto 0);
  signal x8_im_DUT_in : std_logic_vector(31 downto 0);
  signal x9_re_DUT_in : std_logic_vector(31 downto 0);
  signal x9_im_DUT_in : std_logic_vector(31 downto 0);
  signal x10_re_DUT_in : std_logic_vector(31 downto 0);
  signal x10_im_DUT_in : std_logic_vector(31 downto 0);
  signal x11_re_DUT_in : std_logic_vector(31 downto 0);
  signal x11_im_DUT_in : std_logic_vector(31 downto 0);
  signal x12_re_DUT_in : std_logic_vector(31 downto 0);
  signal x12_im_DUT_in : std_logic_vector(31 downto 0);
  signal x13_re_DUT_in : std_logic_vector(31 downto 0);
  signal x13_im_DUT_in : std_logic_vector(31 downto 0);
  signal x14_re_DUT_in : std_logic_vector(31 downto 0);
  signal x14_im_DUT_in : std_logic_vector(31 downto 0);
  signal x15_re_DUT_in : std_logic_vector(31 downto 0);
  signal x15_im_DUT_in : std_logic_vector(31 downto 0);
  signal y0_re_DUT_out : std_logic_vector(31 downto 0);
  signal y0_im_DUT_out : std_logic_vector(31 downto 0);
  signal y1_re_DUT_out : std_logic_vector(31 downto 0);
  signal y1_im_DUT_out : std_logic_vector(31 downto 0);
  signal y2_re_DUT_out : std_logic_vector(31 downto 0);
  signal y2_im_DUT_out : std_logic_vector(31 downto 0);
  signal y3_re_DUT_out : std_logic_vector(31 downto 0);
  signal y3_im_DUT_out : std_logic_vector(31 downto 0);
  signal y4_re_DUT_out : std_logic_vector(31 downto 0);
  signal y4_im_DUT_out : std_logic_vector(31 downto 0);
  signal y5_re_DUT_out : std_logic_vector(31 downto 0);
  signal y5_im_DUT_out : std_logic_vector(31 downto 0);
  signal y6_re_DUT_out : std_logic_vector(31 downto 0);
  signal y6_im_DUT_out : std_logic_vector(31 downto 0);
  signal y7_re_DUT_out : std_logic_vector(31 downto 0);
  signal y7_im_DUT_out : std_logic_vector(31 downto 0);
  signal y8_re_DUT_out : std_logic_vector(31 downto 0);
  signal y8_im_DUT_out : std_logic_vector(31 downto 0);
  signal y9_re_DUT_out : std_logic_vector(31 downto 0);
  signal y9_im_DUT_out : std_logic_vector(31 downto 0);
  signal y10_re_DUT_out : std_logic_vector(31 downto 0);
  signal y10_im_DUT_out : std_logic_vector(31 downto 0);
  signal y11_re_DUT_out : std_logic_vector(31 downto 0);
  signal y11_im_DUT_out : std_logic_vector(31 downto 0);
  signal y12_re_DUT_out : std_logic_vector(31 downto 0);
  signal y12_im_DUT_out : std_logic_vector(31 downto 0);
  signal y13_re_DUT_out : std_logic_vector(31 downto 0);
  signal y13_im_DUT_out : std_logic_vector(31 downto 0);
  signal y14_re_DUT_out : std_logic_vector(31 downto 0);
  signal y14_im_DUT_out : std_logic_vector(31 downto 0);
  signal y15_re_DUT_out : std_logic_vector(31 downto 0);
  signal y15_im_DUT_out : std_logic_vector(31 downto 0);
  type output_mux_input_t is array (0 to 31) of std_logic_vector(31 downto 0);
  signal output_mux_input : output_mux_input_t;

  begin
    DUT : entity work.implementedSystem_toplevel
      port map (
        clk => clk,
        rst => rst,
        x0_re => x0_re_DUT_in,
        x0_im => x0_im_DUT_in,
        x1_re => x1_re_DUT_in,
        x1_im => x1_im_DUT_in,
        x2_re => x2_re_DUT_in,
        x2_im => x2_im_DUT_in,
        x3_re => x3_re_DUT_in,
        x3_im => x3_im_DUT_in,
        x4_re => x4_re_DUT_in,
        x4_im => x4_im_DUT_in,
        x5_re => x5_re_DUT_in,
        x5_im => x5_im_DUT_in,
        x6_re => x6_re_DUT_in,
        x6_im => x6_im_DUT_in,
        x7_re => x7_re_DUT_in,
        x7_im => x7_im_DUT_in,
        x8_re => x8_re_DUT_in,
        x8_im => x8_im_DUT_in,
        x9_re => x9_re_DUT_in,
        x9_im => x9_im_DUT_in,
        x10_re => x10_re_DUT_in,
        x10_im => x10_im_DUT_in,
        x11_re => x11_re_DUT_in,
        x11_im => x11_im_DUT_in,
        x12_re => x12_re_DUT_in,
        x12_im => x12_im_DUT_in,
        x13_re => x13_re_DUT_in,
        x13_im => x13_im_DUT_in,
        x14_re => x14_re_DUT_in,
        x14_im => x14_im_DUT_in,
        x15_re => x15_re_DUT_in,
        x15_im => x15_im_DUT_in,
        y0_re => y0_re_DUT_out,
        y0_im => y0_im_DUT_out,
        y1_re => y1_re_DUT_out,
        y1_im => y1_im_DUT_out,
        y2_re => y2_re_DUT_out,
        y2_im => y2_im_DUT_out,
        y3_re => y3_re_DUT_out,
        y3_im => y3_im_DUT_out,
        y4_re => y4_re_DUT_out,
        y4_im => y4_im_DUT_out,
        y5_re => y5_re_DUT_out,
        y5_im => y5_im_DUT_out,
        y6_re => y6_re_DUT_out,
        y6_im => y6_im_DUT_out,
        y7_re => y7_re_DUT_out,
        y7_im => y7_im_DUT_out,
        y8_re => y8_re_DUT_out,
        y8_im => y8_im_DUT_out,
        y9_re => y9_re_DUT_out,
        y9_im => y9_im_DUT_out,
        y10_re => y10_re_DUT_out,
        y10_im => y10_im_DUT_out,
        y11_re => y11_re_DUT_out,
        y11_im => y11_im_DUT_out,
        y12_re => y12_re_DUT_out,
        y12_im => y12_im_DUT_out,
        y13_re => y13_re_DUT_out,
        y13_im => y13_im_DUT_out,
        y14_re => y14_re_DUT_out,
        y14_im => y14_im_DUT_out,
        y15_re => y15_re_DUT_out,
        y15_im => y15_im_DUT_out
       );
    process(clk)
      begin
        if (rising_edge(clk)) then
          if (x0_re_enable = '1') then
            x0_re_DUT_in <= shared_input;
          end if; -- enable for input x0_re
          if (x0_im_enable = '1') then
            x0_im_DUT_in <= shared_input;
          end if; -- enable for input x0_im
          if (x1_re_enable = '1') then
            x1_re_DUT_in <= shared_input;
          end if; -- enable for input x1_re
          if (x1_im_enable = '1') then
            x1_im_DUT_in <= shared_input;
          end if; -- enable for input x1_im
          if (x2_re_enable = '1') then
            x2_re_DUT_in <= shared_input;
          end if; -- enable for input x2_re
          if (x2_im_enable = '1') then
            x2_im_DUT_in <= shared_input;
          end if; -- enable for input x2_im
          if (x3_re_enable = '1') then
            x3_re_DUT_in <= shared_input;
          end if; -- enable for input x3_re
          if (x3_im_enable = '1') then
            x3_im_DUT_in <= shared_input;
          end if; -- enable for input x3_im
          if (x4_re_enable = '1') then
            x4_re_DUT_in <= shared_input;
          end if; -- enable for input x4_re
          if (x4_im_enable = '1') then
            x4_im_DUT_in <= shared_input;
          end if; -- enable for input x4_im
          if (x5_re_enable = '1') then
            x5_re_DUT_in <= shared_input;
          end if; -- enable for input x5_re
          if (x5_im_enable = '1') then
            x5_im_DUT_in <= shared_input;
          end if; -- enable for input x5_im
          if (x6_re_enable = '1') then
            x6_re_DUT_in <= shared_input;
          end if; -- enable for input x6_re
          if (x6_im_enable = '1') then
            x6_im_DUT_in <= shared_input;
          end if; -- enable for input x6_im
          if (x7_re_enable = '1') then
            x7_re_DUT_in <= shared_input;
          end if; -- enable for input x7_re
          if (x7_im_enable = '1') then
            x7_im_DUT_in <= shared_input;
          end if; -- enable for input x7_im
          if (x8_re_enable = '1') then
            x8_re_DUT_in <= shared_input;
          end if; -- enable for input x8_re
          if (x8_im_enable = '1') then
            x8_im_DUT_in <= shared_input;
          end if; -- enable for input x8_im
          if (x9_re_enable = '1') then
            x9_re_DUT_in <= shared_input;
          end if; -- enable for input x9_re
          if (x9_im_enable = '1') then
            x9_im_DUT_in <= shared_input;
          end if; -- enable for input x9_im
          if (x10_re_enable = '1') then
            x10_re_DUT_in <= shared_input;
          end if; -- enable for input x10_re
          if (x10_im_enable = '1') then
            x10_im_DUT_in <= shared_input;
          end if; -- enable for input x10_im
          if (x11_re_enable = '1') then
            x11_re_DUT_in <= shared_input;
          end if; -- enable for input x11_re
          if (x11_im_enable = '1') then
            x11_im_DUT_in <= shared_input;
          end if; -- enable for input x11_im
          if (x12_re_enable = '1') then
            x12_re_DUT_in <= shared_input;
          end if; -- enable for input x12_re
          if (x12_im_enable = '1') then
            x12_im_DUT_in <= shared_input;
          end if; -- enable for input x12_im
          if (x13_re_enable = '1') then
            x13_re_DUT_in <= shared_input;
          end if; -- enable for input x13_re
          if (x13_im_enable = '1') then
            x13_im_DUT_in <= shared_input;
          end if; -- enable for input x13_im
          if (x14_re_enable = '1') then
            x14_re_DUT_in <= shared_input;
          end if; -- enable for input x14_re
          if (x14_im_enable = '1') then
            x14_im_DUT_in <= shared_input;
          end if; -- enable for input x14_im
          if (x15_re_enable = '1') then
            x15_re_DUT_in <= shared_input;
          end if; -- enable for input x15_re
          if (x15_im_enable = '1') then
            x15_im_DUT_in <= shared_input;
          end if; -- enable for input x15_im
        end if; -- clk
      end process;
    output_mux_input(0) <= y0_re_DUT_out;
    output_mux_input(1) <= y0_im_DUT_out;
    output_mux_input(2) <= y1_re_DUT_out;
    output_mux_input(3) <= y1_im_DUT_out;
    output_mux_input(4) <= y2_re_DUT_out;
    output_mux_input(5) <= y2_im_DUT_out;
    output_mux_input(6) <= y3_re_DUT_out;
    output_mux_input(7) <= y3_im_DUT_out;
    output_mux_input(8) <= y4_re_DUT_out;
    output_mux_input(9) <= y4_im_DUT_out;
    output_mux_input(10) <= y5_re_DUT_out;
    output_mux_input(11) <= y5_im_DUT_out;
    output_mux_input(12) <= y6_re_DUT_out;
    output_mux_input(13) <= y6_im_DUT_out;
    output_mux_input(14) <= y7_re_DUT_out;
    output_mux_input(15) <= y7_im_DUT_out;
    output_mux_input(16) <= y8_re_DUT_out;
    output_mux_input(17) <= y8_im_DUT_out;
    output_mux_input(18) <= y9_re_DUT_out;
    output_mux_input(19) <= y9_im_DUT_out;
    output_mux_input(20) <= y10_re_DUT_out;
    output_mux_input(21) <= y10_im_DUT_out;
    output_mux_input(22) <= y11_re_DUT_out;
    output_mux_input(23) <= y11_im_DUT_out;
    output_mux_input(24) <= y12_re_DUT_out;
    output_mux_input(25) <= y12_im_DUT_out;
    output_mux_input(26) <= y13_re_DUT_out;
    output_mux_input(27) <= y13_im_DUT_out;
    output_mux_input(28) <= y14_re_DUT_out;
    output_mux_input(29) <= y14_im_DUT_out;
    output_mux_input(30) <= y15_re_DUT_out;
    output_mux_input(31) <= y15_im_DUT_out;
    shared_output <= output_mux_input(to_integer(unsigned(output_select)));
    
end architecture;
